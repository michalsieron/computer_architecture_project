`timescale 1ps/1ps

`include "fadd_a1.v"

module fadd_a1_tb;

reg [31:0] a, b;
wire [31:0] out;

reg clk = 1'b1;

fadd_a1 uut(a, b, out);

always clk = #5 ~clk;

initial begin

	$dumpfile("fadd_a1_out.vcd");
	$dumpvars(0, fadd_a1_tb);
	test_case(32'hdfe30df6, 32'h5ec6bdb6);
	test_case(32'h5e53fd68, 32'hdee630bf);
	test_case(32'hdf5b5ce9, 32'h5f5fde8b);
	test_case(32'hdeddc6d9, 32'hde58a76f);
	test_case(32'hdf736e8a, 32'hde677a15);
	test_case(32'h5ec991ed, 32'hdefa2e7f);
	test_case(32'h5efbaefb, 32'hde72f03a);
	test_case(32'h5ff86638, 32'h5fef6580);
	test_case(32'hdedfb03f, 32'h5fd53362);
	test_case(32'hdefc8d25, 32'h5fc8e900);
	test_case(32'h5ff7f1a5, 32'hdf475325);
	test_case(32'hdfdf2602, 32'hdf64beb1);
	test_case(32'hdfcfc3b7, 32'hde7ce839);
	test_case(32'h5ff2b9b8, 32'h5fd78a0d);
	test_case(32'hdfd578dd, 32'h5efb6ab3);
	test_case(32'h5ee25a22, 32'hde73d559);
	test_case(32'hdf4f24b5, 32'h5ecb1b4d);
	test_case(32'hdffbf504, 32'hdfde817d);
	test_case(32'hdf6f1fd7, 32'h5f64e0da);
	test_case(32'h5fc37724, 32'hddf6c139);
	test_case(32'h5fe43b57, 32'hdff5a96d);
	test_case(32'h5ff7c141, 32'hde5943cc);
	test_case(32'hde787c9d, 32'hdfe191a7);
	test_case(32'hdff5c0c9, 32'h5fef67d1);
	test_case(32'h5ff9904a, 32'hde619e45);
	test_case(32'h5fef0246, 32'h5fe019de);
	test_case(32'h5fef37f5, 32'hdee4df58);
	test_case(32'h5fd05d1a, 32'h5cf976eb);
	test_case(32'hdfcf3543, 32'hdfc6769d);
	test_case(32'h5e439733, 32'hdfd2d603);
	test_case(32'h5edbfe3d, 32'h5f591037);
	test_case(32'h5fc67c08, 32'h5ffb9666);
	test_case(32'h5fe6472f, 32'hdfe835f4);
	test_case(32'h5f46fb0a, 32'h5feed653);
	test_case(32'hded1d8d8, 32'h5bc71d03);
	test_case(32'hdffd6c44, 32'h5fd4258f);
	test_case(32'hdf6e8e49, 32'hdecce38f);
	test_case(32'h5fe422d2, 32'h5fc3e2ed);
	test_case(32'hdfed7da6, 32'hdfcce49a);
	test_case(32'h5ff18bb2, 32'hded2ed55);
	test_case(32'h5f4ca068, 32'hdff08db5);
	test_case(32'h5e6262d6, 32'h5f7b3ab1);
	test_case(32'h5ff73559, 32'hdfcd10fa);
	test_case(32'hde505a5c, 32'h5ed5ca4c);
	test_case(32'h5fcd3a79, 32'hdeca8553);
	test_case(32'h5fce4afb, 32'h5d73f667);
	test_case(32'h5f45ed9f, 32'h5fec9c36);
	test_case(32'h5f7a3186, 32'hdf416342);
	test_case(32'hdfda4421, 32'hdd76ea21);
	test_case(32'h5ffa0f48, 32'hdfe5f451);
	test_case(32'hdf591597, 32'hdffd6f2c);
	test_case(32'hdf40810f, 32'h5f638b17);
	test_case(32'h5fd6ff43, 32'h5fcb907f);
	test_case(32'h5fef1c6d, 32'h5f7cec09);
	test_case(32'hdff80fd7, 32'h5ec4ef69);
	test_case(32'hdfeed3a3, 32'h5ff7a0b1);
	test_case(32'hdd743c89, 32'h5fc442e5);
	test_case(32'h5fdff311, 32'h5e76fd10);
	test_case(32'h5fd43231, 32'hdfd31c2d);
	test_case(32'hdec80b17, 32'h5fefe5fc);
	test_case(32'h5e497f02, 32'h5e636529);
	test_case(32'hdfc08171, 32'hdfe29527);
	test_case(32'h5fef123f, 32'h5fd9a87b);
	test_case(32'hdfd9288d, 32'h5ef0fc43);
	test_case(32'hdde7ca75, 32'h5fd9cd1c);
	test_case(32'h5fc8c759, 32'hded72c28);
	test_case(32'hdf658e69, 32'hdfd5a8fb);
	test_case(32'h5ffffa3c, 32'h5fcc89ef);
	test_case(32'h5dc4a2fd, 32'h5fceeabc);
	test_case(32'h5ef086a9, 32'h5cca32ef);
	test_case(32'h5e5ee68f, 32'h5f5a75a5);
	test_case(32'hdfe8afc3, 32'h5f705726);
	test_case(32'h5ff6547b, 32'h5fff459e);
	test_case(32'h5eee07be, 32'hdf771798);
	test_case(32'h5f4ecb1e, 32'h5fec6d45);
	test_case(32'hdfd519b3, 32'h5f7d4e44);
	test_case(32'hdd5d9f80, 32'hde62b9c9);
	test_case(32'h5f7142f3, 32'hdf541031);
	test_case(32'hde4a9dc1, 32'h5f6dcf3c);
	test_case(32'hdfec663c, 32'hdfd7acda);
	test_case(32'h5fe00e5c, 32'h5f4cc403);
	test_case(32'hdfd416e2, 32'h5ffbede0);
	test_case(32'hdfc79fea, 32'h5fe79d43);
	test_case(32'hdfdb34fc, 32'hdefdf92c);
	test_case(32'hdf72ddef, 32'h5fdb7a4d);
	test_case(32'hdfe7950f, 32'h5fcb13a2);
	test_case(32'hdf5192fb, 32'h5f448db7);
	test_case(32'h5ff245b1, 32'h5e7ff623);
	test_case(32'h5ff6c035, 32'hdfd8a17b);
	test_case(32'h5e5d44bf, 32'hde7110fa);
	test_case(32'h5fcbcddf, 32'h5efe8f80);
	test_case(32'h5efb87a1, 32'h5f533a94);
	test_case(32'h5fcaa951, 32'hdff9e95c);
	test_case(32'hdf7b8400, 32'hdf5dd866);
	test_case(32'hdf68e66e, 32'h5fe23209);
	test_case(32'hdf70abff, 32'hdff23c1a);
	test_case(32'hdfc89a79, 32'h5fc1c61b);
	test_case(32'hdfc8b6ca, 32'hdeec950e);
	test_case(32'hdfcae845, 32'hddf317bb);
	test_case(32'hdf79e48e, 32'h5fe15835);
	test_case(32'hdfd9d7cb, 32'h5f770ff7);
	test_case(32'hdefecd6e, 32'hdf649484);
	test_case(32'hdfc60919, 32'hdff72944);
	test_case(32'h5f6401f8, 32'h5f7fa914);
	test_case(32'hdfc2d30b, 32'h5ec0569b);
	test_case(32'h5ff71904, 32'h5f6829c8);
	test_case(32'h5bf32e1f, 32'h5fec039a);
	test_case(32'h5e452a7f, 32'hdec01c4a);
	test_case(32'h5e5c16f6, 32'h5fd1fe2f);
	test_case(32'hdfdffd75, 32'hdfee7adb);
	test_case(32'h5fde3211, 32'hde7b6225);
	test_case(32'hddcbe034, 32'hddf7270e);
	test_case(32'h5fd1ef46, 32'h5fc09bd7);
	test_case(32'h5fd24150, 32'h5fd0d651);
	test_case(32'h5ffcfa32, 32'hde6d95b4);
	test_case(32'hde44f3ac, 32'h5de9df4b);
	test_case(32'hdf4af68f, 32'h5f56656e);
	test_case(32'hdf6e0f33, 32'h5ed72138);
	test_case(32'hdfc9da9c, 32'hde6c7517);
	test_case(32'hdff7e112, 32'h5f5d7b06);
	test_case(32'hdf510f4c, 32'hdfc55234);
	test_case(32'h5edd3c2d, 32'h5fecb912);
	test_case(32'h5fd4bd0a, 32'h5f78bb62);
	test_case(32'h5f42f1a2, 32'hdfc6100d);
	test_case(32'hdfc13ccc, 32'h5f780469);
	test_case(32'h5ffc44f8, 32'h5cee2c50);
	test_case(32'hdfc9f9dc, 32'hdec1245a);
	test_case(32'hdfc1c50e, 32'hdfcd49a8);
	test_case(32'hdee1c03c, 32'hdf7b32fa);
	test_case(32'h5f569317, 32'h5fdde096);
	test_case(32'h5f4e14dc, 32'hde5ff180);
	test_case(32'hded704c9, 32'h5fd8ddbc);
	test_case(32'h5ec2aa61, 32'h5fc1462a);
	test_case(32'h5f70c5da, 32'hdfd359fd);
	test_case(32'h5ffd0cfc, 32'hdfe2fd8c);
	test_case(32'hdfde7c7a, 32'h5ff2de9e);
	test_case(32'h5ff8fb86, 32'hdf73e26b);
	test_case(32'h5ed0932c, 32'hdfc8071a);
	test_case(32'hdf4fe39f, 32'h5eda391c);
	test_case(32'hdef7f40e, 32'h5f6400f2);
	test_case(32'h5e7223e8, 32'h5fc4e5bf);
	test_case(32'h5fea2235, 32'hdfea302f);
	test_case(32'hdf4f0c26, 32'hdfea4d68);
	test_case(32'h5fd96b8c, 32'h5fc9c64b);
	test_case(32'hdffda9f6, 32'hdff21bb6);
	test_case(32'hded14255, 32'h5f6d9628);
	test_case(32'hdfef15ea, 32'hdffd070e);
	test_case(32'hdf7fc0af, 32'hdfc797f8);
	test_case(32'hdfc95b3e, 32'hdf71b619);
	test_case(32'h5e72f36a, 32'h5fcd7486);
	test_case(32'hdf57a4b6, 32'h5e7c4c74);
	test_case(32'hdfffc019, 32'h5feddccd);
	test_case(32'h5e43c754, 32'h5f687236);
	test_case(32'hdf67985d, 32'h5fec4b1d);
	test_case(32'h5f6312fe, 32'h5fc3cb56);
	test_case(32'h5fd4ec7d, 32'h5fe30a05);
	test_case(32'h5ff36eb0, 32'h5e52b753);
	test_case(32'hdf660533, 32'hdfd9686e);
	test_case(32'hdfc2e6f8, 32'h5f755f43);
	test_case(32'h5e6f0add, 32'hde495618);
	test_case(32'hdf45dc03, 32'h5ff066a9);
	test_case(32'h5f4efc87, 32'hdffc4c64);
	test_case(32'hdeec330e, 32'hdecca054);
	test_case(32'h5f4fc0b7, 32'h5f59905f);
	test_case(32'hdecca34f, 32'hdf7852c0);
	test_case(32'h5ef38cba, 32'hdfe6f0c5);
	test_case(32'h5fdc05c1, 32'h5fd0c44f);
	test_case(32'h5f74e8fb, 32'h5efb3518);
	test_case(32'h5ff5554c, 32'h5ed49f6b);
	test_case(32'h5f795d73, 32'hdf5a9192);
	test_case(32'hdf49327b, 32'h5ffee263);
	test_case(32'h5ffae563, 32'hdff12f6b);
	test_case(32'hde753c58, 32'h5fc98341);
	test_case(32'h5fcaf1c9, 32'h5f73b1b5);
	test_case(32'h5ee5f358, 32'h5f781283);
	test_case(32'h5fcecee8, 32'h5feb6a7a);
	test_case(32'hdfdb85c0, 32'h5ffe71aa);
	test_case(32'h5efe2d6f, 32'hdfd52d7f);
	test_case(32'h5c5af798, 32'h5ee4b67e);
	test_case(32'h5fc4e305, 32'hdfca135e);
	test_case(32'h5ec671c3, 32'hdfd81b6e);
	test_case(32'hdf582192, 32'hdffed2d2);
	test_case(32'hdeda99c8, 32'hdf798586);
	test_case(32'h5e530698, 32'hdffe1642);
	test_case(32'hdf770b7c, 32'h5f7e4e1a);
	test_case(32'h5ff2b2c3, 32'hdfe95442);
	test_case(32'hdedd5fb8, 32'hdf767827);
	test_case(32'hdfca81db, 32'hdf4e7e54);
	test_case(32'hdfd3d88a, 32'hdf607051);
	test_case(32'hdfc5e778, 32'hdf660c05);
	test_case(32'h5eeee971, 32'h5e672f38);
	test_case(32'h5fcd595e, 32'hdfe4db05);
	test_case(32'hdf5008eb, 32'hdf69aa1a);
	test_case(32'h5fc66a6a, 32'hdf763702);
	test_case(32'h5fdaf626, 32'hdff5c50e);
	test_case(32'h5ff886e5, 32'h5fe776ef);
	test_case(32'h5f7d1756, 32'h5d4658da);
	test_case(32'hdfd93af7, 32'h5ed4fbd8);
	test_case(32'h5fe565cf, 32'hdfecb816);
	test_case(32'hded54598, 32'h5fd7a8bd);
	test_case(32'h5fdf106c, 32'h5fd1d8d1);
	test_case(32'h5fec2b55, 32'hdce1efca);
	test_case(32'h5e748ddd, 32'h5fce3e2f);
	test_case(32'hdf4e6785, 32'h5fee6e58);
	test_case(32'hdf634c5b, 32'h5f5cbd1f);
	test_case(32'hdfe40941, 32'hdfe1119b);
	test_case(32'h5dc70562, 32'hdfce78fb);
	test_case(32'h5edb919c, 32'h5f5e768b);
	test_case(32'h5fcc882a, 32'h5ffe0f1e);
	test_case(32'h5ee28540, 32'hdfc1ef4a);
	test_case(32'hdfec733a, 32'hdfdf9c80);
	test_case(32'h5e6fac1a, 32'h5a703deb);
	test_case(32'hdfd97fd2, 32'hdffa8258);
	test_case(32'h5f6cd528, 32'hdfdb55fa);
	test_case(32'h5e6bd512, 32'h5ffab524);
	test_case(32'hdfe09197, 32'h5e4202d9);
	test_case(32'hde5709c4, 32'h5e763b10);
	test_case(32'hdedb89fa, 32'h5fff122e);
	test_case(32'hdf416f4e, 32'hde62be47);
	test_case(32'hdff41ae4, 32'h5ef1f4a6);
	test_case(32'h5f458d4a, 32'h5f49d0dd);
	test_case(32'h5f483c4b, 32'h5ee7d5a9);
	test_case(32'hdf46dc94, 32'h5f4197df);
	test_case(32'h5fd1a3b8, 32'h5ff341d1);
	test_case(32'hdf53c5eb, 32'h5fd92bb2);
	test_case(32'h5e5b204d, 32'h5fc3dbef);
	test_case(32'hdf59f1df, 32'h5efa04c5);
	test_case(32'h5ed30445, 32'h5fcaa1a7);
	test_case(32'hdfc28e5d, 32'h5fc37abd);
	test_case(32'h5ec64a04, 32'hdffb027f);
	test_case(32'hdf6a38bf, 32'hddca381d);
	test_case(32'hdfd655cb, 32'hdec3d9b7);
	test_case(32'hdf7e9a6f, 32'h5feac69f);
	test_case(32'h5f774ed1, 32'h5ff21f9a);
	test_case(32'h5fcea059, 32'h5f62eaed);
	test_case(32'hdf5ac7b2, 32'hdf71236d);
	test_case(32'hdff27834, 32'h5ff2b5b1);
	test_case(32'hdf697dd4, 32'hdfd987c7);
	test_case(32'h5fe6c306, 32'hdfcb2c91);
	test_case(32'hdfee436b, 32'hdffb0e53);
	test_case(32'hdfcc31c7, 32'h5feab558);
	test_case(32'h5dd1e357, 32'hde7c1e01);
	test_case(32'hdf6e8249, 32'hdfe42ff6);
	test_case(32'h5fd616fc, 32'h5ffa2aa4);
	test_case(32'h5fecd372, 32'hdff042e1);
	test_case(32'hdf54e5bc, 32'hdf729c8e);
	test_case(32'hded018f0, 32'hdfef35a2);
	test_case(32'h5e485f7e, 32'hdf47996f);
	test_case(32'hdfd524f0, 32'hdfc5dd37);
	test_case(32'hdffb0838, 32'h5fcd50e9);
	test_case(32'hdfdd8a26, 32'h5fc95383);
	test_case(32'h5fd4fc13, 32'hdfc08754);
	test_case(32'hdedf9fe6, 32'hdfdc875d);
	test_case(32'h5ec69623, 32'hdffb4509);
	test_case(32'hdf467b97, 32'h5ff2bdde);
	test_case(32'h5f65a867, 32'h5fc678f7);
	test_case(32'hdfd69c0b, 32'hddc6c928);
	test_case(32'h5e7c57d4, 32'h5ef22a8b);
	test_case(32'h5eca3e08, 32'hdf46e22f);
	test_case(32'h5fee4d33, 32'hdfc31a2f);
	test_case(32'hddc232a8, 32'h5fc776bc);
	test_case(32'h5e7eb475, 32'hdf6df3d8);
	test_case(32'hdfc8ad72, 32'h5f638e0d);
	test_case(32'h5eee4d8e, 32'hdfe8dd5f);
	test_case(32'hdff2351e, 32'hdfc996ee);
	test_case(32'hdd56c0ed, 32'hdfec524d);
	test_case(32'hdfd922ac, 32'hdfee9036);
	test_case(32'h5e5226c1, 32'h5fe1152a);
	test_case(32'hdf5e8f9f, 32'hdf673b8c);
	test_case(32'h5ff2e6d0, 32'h5d5abd67);
	test_case(32'hdf44bac3, 32'h5edf1071);
	test_case(32'hdffdf5d1, 32'h5f763e4e);
	test_case(32'hdfe3abfd, 32'hdfe87d5b);
	test_case(32'h5f6631a5, 32'hdf542eb6);
	test_case(32'h5ef8510d, 32'hdfcb4ba9);
	test_case(32'hdfcb5546, 32'h5e5bd37f);
	test_case(32'hdffab6a3, 32'hdff8f7e2);
	test_case(32'h5ff62fe6, 32'hdf7d9ccb);
	test_case(32'h5f4f0d3c, 32'h5fc21977);
	test_case(32'h5afd6647, 32'hdff0e2b5);
	test_case(32'h5fff0273, 32'hdfc2cba4);
	test_case(32'hdff63eaa, 32'h5fd5f7d2);
	test_case(32'h5f58363e, 32'h5f43f7f9);
	test_case(32'h5fc79c39, 32'h5fe67f12);
	test_case(32'h5fe33dbc, 32'hdfe97a36);
	test_case(32'h5ff990cc, 32'h5ffa66d3);
	test_case(32'hdf4ed43d, 32'h5edde82e);
	test_case(32'h5dd02a25, 32'hdde39c49);
	test_case(32'hddfa5471, 32'hdff01b67);
	test_case(32'h5ed41b8b, 32'hdfe51a62);
	test_case(32'hdfc7c2da, 32'hdf52a3a2);
	test_case(32'h5ed37852, 32'hdefc9e7f);
	test_case(32'h5fc99f72, 32'h5f479c03);
	test_case(32'hdf707744, 32'hdf4137b7);
	test_case(32'h5cffcf78, 32'h5fc5509c);
	test_case(32'h5e69d8e5, 32'hdee511b4);
	test_case(32'h5e407798, 32'hdfc50edc);
	test_case(32'h5ffec5fb, 32'h5ff432f7);
	test_case(32'h5ede903c, 32'hdedb1c7e);
	test_case(32'h5ff2350d, 32'hddc1b19d);
	test_case(32'hdfc0bce6, 32'hdf4c68cc);
	test_case(32'h5fec6e87, 32'h5f6bf7d8);
	test_case(32'h5fcb50d7, 32'hdfdef204);
	test_case(32'hdffdbd09, 32'hdee94668);
	test_case(32'h5f69b3b7, 32'hdfdf6ae8);
	test_case(32'h5feda093, 32'hdfde8ea4);
	test_case(32'h5d482ae7, 32'h5fc8d9cc);
	test_case(32'hdfd01e76, 32'hdfee7a92);
	test_case(32'h5e5eb5ae, 32'h5f5d4292);
	test_case(32'hdde4616e, 32'h5fd90dcc);
	test_case(32'h5fda041d, 32'h5ff2fae7);
	test_case(32'h5f4ab9f5, 32'hdec78415);
	test_case(32'h5eeb4908, 32'h5fd4f7c0);
	test_case(32'hdfe80157, 32'h5fed7adf);
	test_case(32'hdfc3a35a, 32'hde64dac6);
	test_case(32'h5f5603ec, 32'h5f7dbe8f);
	test_case(32'h5d5b180d, 32'h5fece746);
	test_case(32'hdf713b0a, 32'h5f6308a4);
	test_case(32'hdfc1df74, 32'hdfc7788a);
	test_case(32'hdfc99da9, 32'h5fcd7f64);
	test_case(32'h5f660d65, 32'h5f77d510);
	test_case(32'hdfdf5f96, 32'hdee55c68);
	test_case(32'h5f4cfb1a, 32'h5feff7aa);
	test_case(32'h5e65abbc, 32'hdfd9e7f1);
	test_case(32'hdf6535c1, 32'hdecc4fca);
	test_case(32'hddd4c9e8, 32'h5de7642e);
	test_case(32'hdf720f7e, 32'h5fe16c25);
	test_case(32'hdf7453d5, 32'h5fd72158);
	test_case(32'hdfef3290, 32'hdf5dddea);
	test_case(32'hdfcc56f2, 32'hdf53c34f);
	test_case(32'h5ed496da, 32'hdecfb8d1);
	test_case(32'h5f79da18, 32'h5f6c8769);
	test_case(32'h5f4795ff, 32'h5fef3a7e);
	test_case(32'hdf764ea3, 32'hdffbc8ae);
	test_case(32'hdf526972, 32'hde4b7370);
	test_case(32'hdeee2a74, 32'h5f578e35);
	test_case(32'h5fc3f2f3, 32'hdff73cfb);
	test_case(32'h5fe75b60, 32'h5fd8140d);
	test_case(32'h5d458486, 32'h5fcb8f07);
	test_case(32'hdfece342, 32'h5fd65bc6);
	test_case(32'hdf5a7ee5, 32'hde43c589);
	test_case(32'h5ffa9bd9, 32'hdefa57dc);
	test_case(32'hdfd4a1a2, 32'hdf647012);
	test_case(32'hdfd209b9, 32'h5f7eb9b0);
	test_case(32'hdd694afd, 32'hdfe64eb9);
	test_case(32'h5ff10060, 32'h5fead3d6);
	test_case(32'hde66269f, 32'h5f43b383);
	test_case(32'h5fc13d6c, 32'h5f6baa74);
	test_case(32'hdffd3ae4, 32'hdf478e6e);
	test_case(32'hdff89f11, 32'h5fe2fbb0);
	test_case(32'h5fe50a34, 32'hdff89f5a);
	test_case(32'h5fde1ca6, 32'hdfd946d8);
	test_case(32'h5fc2bdcf, 32'h5ff90967);
	test_case(32'h5fde79cd, 32'hdfd5d254);
	test_case(32'h5fd8ea1a, 32'hdee56103);
	test_case(32'hdff0f1ab, 32'hdf4c1467);
	test_case(32'hdf770782, 32'hdff4d9ca);
	test_case(32'hdf76d1a0, 32'h5f74598f);
	test_case(32'h5fd928a5, 32'h5fd7f0b5);
	test_case(32'h5fe9e099, 32'hdff86884);
	test_case(32'hde7a5c06, 32'hdfe46130);
	test_case(32'h5ef1f47a, 32'h5fe781fa);
	test_case(32'h5f761625, 32'h5ff9a6fa);
	test_case(32'h5ec6f358, 32'hdfd7b623);
	test_case(32'h5ff56d07, 32'hdeda3158);
	test_case(32'h5f6ee701, 32'hdf5fffd5);
	test_case(32'hdf6826e9, 32'hdf5c7c11);
	test_case(32'hdff85f66, 32'hdffe785d);
	test_case(32'hdfd356b5, 32'hdfde6a74);
	test_case(32'hdfd7b3c4, 32'hdcd46788);
	test_case(32'hdf402f77, 32'hdfc50e60);
	test_case(32'h5ffa7d88, 32'h5f7d6ddb);
	test_case(32'hdee13084, 32'hde778037);
	test_case(32'hde683c85, 32'h5fd8a530);
	test_case(32'hdfee82a5, 32'h5fd3b9d0);
	test_case(32'hdfe9e23b, 32'h5fd528bd);
	test_case(32'h5dde74cf, 32'hdfe40af2);
	test_case(32'h5f5417ee, 32'h5fd77cae);
	test_case(32'hdf7793fb, 32'hdfd06c9c);
	test_case(32'h5f58e657, 32'hdfe21f2c);
	test_case(32'h5fc4e00b, 32'hdfdba06d);
	test_case(32'h5ff756d7, 32'h5ec9eea0);
	test_case(32'h5fe93b37, 32'h5fc2aa44);
	test_case(32'hdedd9704, 32'h5f54e264);
	test_case(32'h5fd9ac64, 32'h5fce307a);
	test_case(32'h5ff7c96b, 32'h5fdf8d95);
	test_case(32'h5fc94916, 32'hdf494693);
	test_case(32'hdf6f2ba5, 32'h5fd1be42);
	test_case(32'h5fd2010d, 32'h5e6a3ca8);
	test_case(32'hdfefdeca, 32'hdf5983ef);
	test_case(32'hdfe1f9d0, 32'h5ece9e05);
	test_case(32'hdfcf5232, 32'hdf6d229f);
	test_case(32'h5f4d89cd, 32'hdfc36cc1);
	test_case(32'h5f63a2a4, 32'hdfccbcb3);
	test_case(32'hdfed0fb1, 32'h5fcfd0f0);
	test_case(32'hdfe46138, 32'h5f6b4f22);
	test_case(32'h5eca74e6, 32'h5ee2b920);
	test_case(32'h5f5edd7e, 32'h5f46a6bc);
	test_case(32'h5fcd044c, 32'h5fcd06a2);
	test_case(32'hdff130b4, 32'hdf5e4908);
	test_case(32'hdff521a3, 32'h5fe8b2db);
	test_case(32'hdfc2ce26, 32'h5ef9e4ec);
	test_case(32'h5fcf8f01, 32'h5feeb1cf);
	test_case(32'h5fd8b220, 32'h5f685524);
	test_case(32'hdf5ca740, 32'h5f4d3fc5);
	test_case(32'h5fce0c25, 32'hdefae971);
	test_case(32'h5f4ae498, 32'hdfe9d8d4);
	test_case(32'h5e780731, 32'h5fe4e0c7);
	test_case(32'h5f70c025, 32'h5fe0d049);
	test_case(32'hdf43023a, 32'h5fef77de);
	test_case(32'h5fd63c72, 32'hdf7710a6);
	test_case(32'h5fd2883c, 32'h5fe7111e);
	test_case(32'hde6a55be, 32'hde619b39);
	test_case(32'hdff886ee, 32'h5fd38000);
	test_case(32'hdefba71c, 32'hdf56f7f7);
	test_case(32'hdfd60ede, 32'hdfda486e);
	test_case(32'hdfc0c523, 32'h5dd5c5b6);
	test_case(32'h5fcaac25, 32'h5fdac8da);
	test_case(32'h5e4eb80d, 32'h5ff92341);
	test_case(32'hdfc70c46, 32'h5c6658b1);
	test_case(32'h5f7733a8, 32'hdfecf1c1);
	test_case(32'hdf411088, 32'hdfdb5024);
	test_case(32'hdf7630f8, 32'h5dd593ac);
	test_case(32'h5f503c77, 32'h5e481a1f);
	test_case(32'h5ed26921, 32'hdef28383);
	test_case(32'hdfc301d0, 32'h5fe73e86);
	test_case(32'h5ee0407c, 32'h5ff5023a);
	test_case(32'h5fc5c776, 32'hdfe7c02c);
	test_case(32'h5fc9a163, 32'hdffd8efc);
	test_case(32'hdfd2ec13, 32'h5ed01247);
	test_case(32'h5fdc3d0e, 32'hdfeb3c7c);
	test_case(32'h5ff57eb2, 32'h5ede6ffe);
	test_case(32'hdfd8d1fe, 32'h5ff767b5);
	test_case(32'h5fef2468, 32'hddd2e3c5);
	test_case(32'h5fef9878, 32'h5d7237a7);
	test_case(32'h5eda6aad, 32'h5feafe47);
	test_case(32'h5f755d58, 32'hdfe8a61e);
	test_case(32'hde537011, 32'h5f6c547e);
	test_case(32'hdf4cdb84, 32'hdfd848b7);
	test_case(32'h5fc1ae87, 32'hded1135a);
	test_case(32'hdfed768d, 32'hdf736680);
	test_case(32'hdfc2632f, 32'h5eec1f47);
	test_case(32'hdf5c62b6, 32'h5e764ea0);
	test_case(32'hdff53452, 32'hdf615608);
	test_case(32'hdfd1456e, 32'h5fdbb3be);
	test_case(32'hdfd5d661, 32'h5e564e47);
	test_case(32'h5e65ffd0, 32'h5ed3bde4);
	test_case(32'h5fd3884e, 32'h5ffdc893);
	test_case(32'h5e637cb6, 32'h5ff031fe);
	test_case(32'hdfc9b3b5, 32'hdf5685c5);
	test_case(32'hde7271e3, 32'hdfd81a8f);
	test_case(32'hdf483ba3, 32'h5f4985c3);
	test_case(32'hdce45ba2, 32'hdd7c6015);
	test_case(32'h5ec14ab6, 32'h5ff36e98);
	test_case(32'h5ecc1111, 32'hdec5a480);
	test_case(32'hdf51e7fa, 32'hdfddb86c);
	test_case(32'h5f437292, 32'hdde98a4a);
	test_case(32'h5f598abf, 32'hdfcafb5b);
	test_case(32'h5f668721, 32'h5e72ae87);
	test_case(32'hdfd96d54, 32'h5fcc1ce5);
	test_case(32'h5ff33021, 32'h5fdf4a36);
	test_case(32'hdff23f5c, 32'hdeec4c7d);
	test_case(32'h5fcbd986, 32'hdfe2e8ae);
	test_case(32'hdee54546, 32'hdf57f1ad);
	test_case(32'hdff2100e, 32'h5f4bd7bb);
	test_case(32'hdfeef39c, 32'h5e75ea8d);
	test_case(32'h5fc774bd, 32'h5fde1b1d);
	test_case(32'hdf6b5006, 32'hdfe120a1);
	test_case(32'hdfd7c8f4, 32'h5e494ff6);
	test_case(32'hdf65fcbe, 32'h5f484e3e);
	test_case(32'h5fd0a03b, 32'h5e410860);
	test_case(32'h5f6f9f31, 32'h5fcca41b);
	test_case(32'hdfe66808, 32'hdfcff3c7);
	test_case(32'h5ff1d378, 32'h5fd9de48);
	test_case(32'hdeca6c19, 32'h5fd3f91c);
	test_case(32'h5f731b6e, 32'hdfcadb55);
	test_case(32'h5ff61e41, 32'h5f538f98);
	test_case(32'hdf784b58, 32'hdf4a94ed);
	test_case(32'h5f451116, 32'h5ff890d1);
	test_case(32'h5f50f0c8, 32'h5ef25f8b);
	test_case(32'hdfdc3e7d, 32'h5fdbe7c4);
	test_case(32'h5fce3082, 32'hdfcbef8b);
	test_case(32'h5f41dbe3, 32'hdf41d828);
	test_case(32'hdf7858d8, 32'hdefc61b1);
	test_case(32'h5fc12aa7, 32'hddd65a98);
	test_case(32'h5f59d8b3, 32'h5ffa2706);
	test_case(32'hdfd3d1df, 32'hdf62a97c);
	test_case(32'hdfd83dfa, 32'h5fed1d26);
	test_case(32'hdef25292, 32'h5fe055e5);
	test_case(32'h5f5d8b2d, 32'hde68f736);
	test_case(32'h5f6881a4, 32'h5fd09633);
	test_case(32'hdfe44413, 32'hdfc196af);
	test_case(32'h5fc79ce5, 32'hdef97eb5);
	test_case(32'h5fe4b2a3, 32'hdde37650);
	test_case(32'h5fd63ce3, 32'h5fea456d);
	test_case(32'h5f4f6721, 32'hdfc48e6a);
	test_case(32'hdfc5f6db, 32'h5fe57175);
	test_case(32'h5f4a1615, 32'h5fef5ab3);
	test_case(32'hdfc3ee50, 32'h5fda4466);
	test_case(32'hdf473346, 32'h5ee1de27);
	test_case(32'h5ecb068b, 32'h5fff56f5);
	test_case(32'hdfec6c39, 32'hde74f09d);
	test_case(32'hdd7bad40, 32'hdff1a518);
	test_case(32'h5e5d4060, 32'hdef53af8);
	test_case(32'h5ffd1b7a, 32'hdf4582cd);
	test_case(32'hdf730f86, 32'hddeca7ca);
	test_case(32'h5fcb5570, 32'h5f6d82cd);
	test_case(32'h5ff5924a, 32'hdfca9999);
	test_case(32'h5d4412bf, 32'h5fd27975);
	test_case(32'h5ff2ae2d, 32'h5fff37de);
	test_case(32'h5fc01ca5, 32'hdee96248);
	test_case(32'h5fc13bb3, 32'h5fcc2cdb);
	test_case(32'hdec6745c, 32'hdffeb8ad);
	test_case(32'h5ed0937c, 32'h5ed2b153);
	test_case(32'h5ec5286d, 32'h5fe6e466);
	test_case(32'hddf7f27a, 32'hdffb2da9);
	test_case(32'hddd7826f, 32'h5dfefd76);
	test_case(32'h5fc0a341, 32'h5e7fb570);
	test_case(32'hdfcd9762, 32'hdfdea1fd);
	test_case(32'hdecf4816, 32'h5f7ec69d);
	test_case(32'h5f686210, 32'hdffc006b);
	test_case(32'hdfcea23a, 32'h5cd7ad99);
	test_case(32'hde77c065, 32'h5f6c1fd6);
	test_case(32'h5fd3e380, 32'h5ffd7f3d);
	test_case(32'hdfd86a3a, 32'h5fc09cd8);
	test_case(32'h5fdd1285, 32'h5fe51c18);
	test_case(32'h5f43aaff, 32'hdf5c8977);
	test_case(32'h5f5332b2, 32'hdec42aaa);
	test_case(32'h5ed9879a, 32'h5ff5b930);
	test_case(32'hdff68c7a, 32'h5ec5abfa);
	test_case(32'hde779e93, 32'h5f5752d9);
	test_case(32'hdffa675c, 32'h5e5675a8);
	test_case(32'h5fce5b50, 32'hdfc1d1c7);
	test_case(32'hdfefb0f8, 32'hdfd81cbf);
	test_case(32'hdfcba1f6, 32'h5fcab9be);
	test_case(32'h5ded5044, 32'h5e7fd5bd);
	test_case(32'hdf4f6139, 32'hdff6eee8);
	test_case(32'h5fc75d7f, 32'hdfc8e0d1);
	test_case(32'h5de366e9, 32'hdffa37ca);
	test_case(32'h5cc77ec2, 32'hdef3b285);
	test_case(32'h5fc2a196, 32'hdf64c02d);
	test_case(32'h5f6bc3aa, 32'hdee93439);
	test_case(32'h5fc0ea3f, 32'hdfc8e983);
	test_case(32'h5fe3dfee, 32'h5f6ad85a);
	test_case(32'h5f64e537, 32'hdfcaf9a0);
	test_case(32'h5ffc7e4e, 32'hdf6481cb);
	test_case(32'hdfc735ac, 32'hdfd21a72);
	test_case(32'hdfc85978, 32'hdf421e29);
	test_case(32'hdfde3d91, 32'h5fddab22);
	test_case(32'hdec2cd07, 32'hded535c9);
	test_case(32'h5feb5909, 32'hdeed85b7);
	test_case(32'h5e54f4a2, 32'h5edf4b3e);
	test_case(32'h5ffd38b2, 32'h5fe36ec9);
	test_case(32'h5f7c0306, 32'hdfd12069);
	test_case(32'h5fcff145, 32'hdff10c90);
	test_case(32'h5fea9a3d, 32'h5fdbc31b);
	test_case(32'h5c7b4f5c, 32'h5def6593);
	test_case(32'hdf67975e, 32'h5fce2146);
	test_case(32'h5fc871fb, 32'hdac24296);
	test_case(32'h5f5d8928, 32'hdfcda43f);
	test_case(32'h5feee857, 32'hdf415f5a);
	test_case(32'h5ee20fef, 32'h5ff8d671);
	test_case(32'h5ec95d1c, 32'hdd4daecd);
	test_case(32'h5ecd1e20, 32'hdfd6acb5);
	test_case(32'h5f4dbae9, 32'h5ff3ba6e);
	test_case(32'hde6ea464, 32'hdfc510a0);
	test_case(32'h5fc636b1, 32'h5fedbcba);
	test_case(32'hdf60d2ec, 32'h5fdb6ffd);
	test_case(32'hdffe0eb0, 32'hdfc42446);
	test_case(32'hdff931d3, 32'h5edb758e);
	test_case(32'hdffb0951, 32'h5fdadc5a);
	test_case(32'h5f5dc2e9, 32'hdfdf8f77);
	test_case(32'h5f57b7ed, 32'hdeeea7e6);
	test_case(32'h5f468bcb, 32'h5f7d7089);
	test_case(32'h5f7bea51, 32'h5e48365b);
	test_case(32'hdfde563f, 32'h5ff8f32b);
	test_case(32'h5dfde7f9, 32'h5d6f6f72);
	test_case(32'hdfc7ace1, 32'h5fdf9848);
	test_case(32'h5fd26ae4, 32'hdfc607a5);
	test_case(32'hdf4c7339, 32'hddcd7292);
	test_case(32'hdf674e1b, 32'hdf66a0da);
	test_case(32'h5fd70712, 32'hdfd4ef0e);
	test_case(32'h5f6d7fd6, 32'h5fdba802);
	test_case(32'hded5da73, 32'h5f75635f);
	test_case(32'h5fc654f9, 32'hdfc948b6);
	test_case(32'hdfc8cae3, 32'hded60d01);
	test_case(32'h5ffe60c5, 32'hde70b640);
	test_case(32'h5fff555e, 32'h5f613d82);
	test_case(32'hdfe17c8f, 32'h5fcdf445);
	test_case(32'h5ff04b76, 32'h5fe783a8);
	test_case(32'hdf565394, 32'h5f4f6872);
	test_case(32'hdfe20be0, 32'hdfc09895);
	test_case(32'h5fcb2c84, 32'h5feb7afa);
	test_case(32'hdfe46bdc, 32'hde747d99);
	test_case(32'hdfcb5837, 32'h5ff6cc58);
	test_case(32'h5ec6930c, 32'hdfcf669e);
	test_case(32'hdfe0e174, 32'h5fec528a);
	test_case(32'hde56122e, 32'h5fda1149);
	test_case(32'h5f5538fd, 32'hdfcc25b5);
	test_case(32'h5fc8f742, 32'h5f4a5453);
	test_case(32'h5fdecb97, 32'hdff0265a);
	test_case(32'hdef76e1d, 32'h5eea9ab3);
	test_case(32'hddeb3338, 32'hdf6d2c8b);
	test_case(32'h5f578dcd, 32'h5fc3a051);
	test_case(32'hdff140fd, 32'h5fe915d5);
	test_case(32'hdfddacf2, 32'h5efc3ee0);
	test_case(32'hdfd6081b, 32'h5ffd8174);
	test_case(32'h5fcc9499, 32'hdfd0be47);
	test_case(32'hdfd02fb3, 32'hdf5966e9);
	test_case(32'h5dff75f1, 32'h5ffce388);
	test_case(32'hdfec3c85, 32'h5df3716a);
	test_case(32'hdfcee61d, 32'hdef9185b);
	test_case(32'h5ff94f96, 32'hde658cf1);
	test_case(32'h5f5d59dd, 32'hdfc3e6c2);
	test_case(32'h5fec41db, 32'hdf744a3b);
	test_case(32'h5fcfa012, 32'hdf66c9a9);
	test_case(32'h5ff736c8, 32'hdde24e75);
	test_case(32'hdf5c69fb, 32'h5f51bb63);
	test_case(32'h5fdfd8ca, 32'hdf7e6ef2);
	test_case(32'h5eecefd6, 32'h5fc93bd9);
	test_case(32'hdfc43b76, 32'h5fe32b67);
	test_case(32'hdf670fec, 32'hdf7c7ba3);
	test_case(32'hdfcd1a4a, 32'h5dfdd900);
	test_case(32'h5fc77f32, 32'h5fceceb2);
	test_case(32'hdf70a7f8, 32'h5edff73c);
	test_case(32'h5f59f773, 32'h5ef8d9f0);
	test_case(32'h5fc6bbdb, 32'hdfc67c6a);
	test_case(32'h5efa9e6c, 32'hdfed593e);
	test_case(32'h5f44664c, 32'hdfeb65bc);
	test_case(32'h5fc76d2e, 32'h5f51259f);
	test_case(32'h5ecaf70d, 32'h5fd9c390);
	test_case(32'hdeca35c9, 32'h5f5d513b);
	test_case(32'h5ff0cc50, 32'h5fe8b0c1);
	test_case(32'h5de84bfa, 32'h5e54f366);
	test_case(32'hdefcd06d, 32'hdf6db3d4);
	test_case(32'hdfc85fe7, 32'hdfefda43);
	test_case(32'h5fd0bfb4, 32'hdffdc18f);
	test_case(32'h5fe2617a, 32'hdfc73fe8);
	test_case(32'h5fd7a2cc, 32'hdf59a9b5);
	test_case(32'hdf657f2a, 32'hdfd27220);
	test_case(32'hded7e1c6, 32'h5f403701);
	test_case(32'h5f424f58, 32'h5fc1e1c2);
	test_case(32'h5e7aa268, 32'h5fcb0a7f);
	test_case(32'h5f5cc004, 32'h5fe413fe);
	test_case(32'h5f4f1dfb, 32'hdf5f5a67);
	test_case(32'hdfc1f93d, 32'hdff66a87);
	test_case(32'hdfc4cf70, 32'hdf77c9ca);
	test_case(32'hdff1bbf5, 32'hdf67619a);
	test_case(32'h5f5e7c62, 32'hdece3532);
	test_case(32'h5fe367ba, 32'hde5f22be);
	test_case(32'h5f6657ea, 32'h5efb1c23);
	test_case(32'h5fed4aa7, 32'hdd5b2bd0);
	test_case(32'h5d7299dd, 32'hdff32ac5);
	test_case(32'h5f41047a, 32'hdfe1344a);
	test_case(32'h5ff0c272, 32'hdff0df80);
	test_case(32'hdffbf8ab, 32'hdfede1ce);
	test_case(32'h5de91c35, 32'h5fea7738);
	test_case(32'h5f78411c, 32'hdffef247);
	test_case(32'h5ff577c1, 32'hdf7828a5);
	test_case(32'hdfcecab1, 32'h5f7e1cc4);
	test_case(32'hdec0466a, 32'h5efa505c);
	test_case(32'hdffa63ba, 32'hdfe31644);
	test_case(32'hde64004c, 32'hdefa36c5);
	test_case(32'h5fe0d267, 32'hdf6c8c42);
	test_case(32'hdfc385a1, 32'hdfc5ea3b);
	test_case(32'hdf6518dd, 32'h5e4d8342);
	test_case(32'h5fe802ee, 32'hdf4a7bbe);
	test_case(32'h5f59a329, 32'h5e6a80ee);
	test_case(32'h5f54698d, 32'h5ffa7d38);
	test_case(32'hde57e362, 32'hdf7d8176);
	test_case(32'hdf45bbd3, 32'hdf4f7a9e);
	test_case(32'h5f612738, 32'hdfedc7aa);
	test_case(32'h5fd9a6e1, 32'hdf40ebb3);
	test_case(32'hdf6e1c0e, 32'h5eeeeb2e);
	test_case(32'hdff3deca, 32'hdfe0f8c3);
	test_case(32'h5f721232, 32'hdf5e7b90);
	test_case(32'hdfc09486, 32'h5fd1de71);
	test_case(32'h5f644af4, 32'hdf75101c);
	test_case(32'h5fc0518c, 32'h5eec46b8);
	test_case(32'hdfc53b51, 32'hdfe89f67);
	test_case(32'h5eef1e1f, 32'hde7f597a);
	test_case(32'hdfcf5abe, 32'hdf5893e6);
	test_case(32'hdfd453e7, 32'hdf4c3a7c);
	test_case(32'h5ffa91d2, 32'hdff06423);
	test_case(32'h5ee933ac, 32'h5feafcec);
	test_case(32'hdd4f65fd, 32'hdf410a6d);
	test_case(32'h5fde8851, 32'hdfc9b09a);
	test_case(32'hdfe50cb3, 32'hdffdfd36);
	test_case(32'h5ece6a09, 32'hdfc33041);
	test_case(32'hdf45d09f, 32'h5ffb40ea);
	test_case(32'hdeceb3a4, 32'hdf5f8072);
	test_case(32'h5ec21bdc, 32'h5ff3aa39);
	test_case(32'h5fc8804d, 32'h5df8876c);
	test_case(32'hdf64b4bc, 32'h5ffac2c9);
	test_case(32'hdeddfce2, 32'hdfd27f15);
	test_case(32'hdfc29758, 32'hdf446ef0);
	test_case(32'hdf64330b, 32'h5fee5b55);
	test_case(32'h5ed03839, 32'h5ee38d9b);
	test_case(32'hdf5e1c97, 32'hdde93666);
	test_case(32'h5fffd690, 32'hdfcd8345);
	test_case(32'hde7db583, 32'hdd718879);
	test_case(32'h5e7f2e9a, 32'h5fd5f290);
	test_case(32'hdfee5dff, 32'h5f51de22);
	test_case(32'h5f5032a0, 32'hdf7ce4fb);
	test_case(32'hdf440f77, 32'h5f5f4659);
	test_case(32'hdf6e09ad, 32'hdf72c1b9);
	test_case(32'h5fddfc91, 32'h5fcbda66);
	test_case(32'hdfdc3cc6, 32'h5fd2e42e);
	test_case(32'h5fdefc9c, 32'hdd663dc6);
	test_case(32'hdfe007cb, 32'hdfdd38a8);
	test_case(32'h5f5222e5, 32'hdf4f6620);
	test_case(32'h5ff7c353, 32'hdee366fe);
	test_case(32'hde61aee8, 32'h5f799751);
	test_case(32'hdf7c74d4, 32'h5e7c78d1);
	test_case(32'hdf5bd1e0, 32'h5f44049a);
	test_case(32'h5f661d10, 32'h5ffac3a8);
	test_case(32'h5fe8766c, 32'hdfea43e8);
	test_case(32'h5f493c53, 32'hdfc3d332);
	test_case(32'hdedb050a, 32'hdfcd4210);
	test_case(32'h5f601483, 32'hdf4623be);
	test_case(32'h5ff9bbe4, 32'hded2189b);
	test_case(32'h5fff37ef, 32'hdeceaaad);
	test_case(32'h5dd200a4, 32'hdff418d8);
	test_case(32'hdffbf8ce, 32'h5ff599d7);
	test_case(32'h5fe93960, 32'h5fff6c96);
	test_case(32'h5fc849cc, 32'h5fd16e99);
	test_case(32'hdf706b28, 32'hdec61dcc);
	test_case(32'hdf66ebdd, 32'hdff7a3b2);
	test_case(32'hdf69a034, 32'hdf709ebe);
	test_case(32'hdfc10233, 32'hde4a0e24);
	test_case(32'hdfc943f0, 32'h5f751235);
	test_case(32'hdff06355, 32'h5ffa473f);
	test_case(32'h5fffdfb0, 32'hdeceaf26);
	test_case(32'h5fc5fb6d, 32'hdfca6207);
	test_case(32'hde56dbcd, 32'h5f7b59d6);
	test_case(32'h5f434500, 32'hdfead2d9);
	test_case(32'h5ff18194, 32'h5fdf547e);
	test_case(32'h5fd54a02, 32'h5eca04eb);
	test_case(32'hdf586984, 32'h5fd125af);
	test_case(32'hdf4c1f93, 32'h5fcf485a);
	test_case(32'h5f68f3f1, 32'hdffe12ee);
	test_case(32'hde52d6f6, 32'h5fd1f661);
	test_case(32'h5fc4134c, 32'hdfc73b0c);
	test_case(32'hdfea15e4, 32'h5eef5b6f);
	test_case(32'hdfd4e2fe, 32'hdf60ec58);
	test_case(32'h5feade3a, 32'hde6b6040);
	test_case(32'h5f513940, 32'hdedabb07);
	test_case(32'hdff71ca0, 32'hde500748);
	test_case(32'hdff23f53, 32'hdfdf6503);
	test_case(32'h5e790252, 32'hde421bf6);
	test_case(32'hdece961e, 32'hdfebb9d8);
	test_case(32'h5ed88292, 32'hdec5380e);
	test_case(32'hdfc08569, 32'h5ed2a5cf);
	test_case(32'h5f623521, 32'hdfff4212);
	test_case(32'hdf5bda49, 32'hdf6a8a01);
	test_case(32'h5c455820, 32'hdfd4fb27);
	test_case(32'h5f76d031, 32'hdd5886d1);
	test_case(32'h5fea01c5, 32'h5fd30b8c);
	test_case(32'h5ff75226, 32'hddc16709);
	test_case(32'hdfd539e5, 32'hdfc72dc5);
	test_case(32'hdff0c6c5, 32'hde4dbf19);
	test_case(32'h5ed7d329, 32'h5ecdf611);
	test_case(32'hde4d3018, 32'hdfdfb2f8);
	test_case(32'hdf4d1fdd, 32'h5fc7ffdd);
	test_case(32'hdf64c3de, 32'h5fca69ce);
	test_case(32'hdee27f91, 32'hdff51b51);
	test_case(32'h5fef8b3f, 32'hdfe1057f);
	test_case(32'hdf4a1aca, 32'hdefa0398);
	test_case(32'hdfec1d43, 32'h5ef93bb6);
	test_case(32'h5ecfbceb, 32'hdfcc74a4);
	test_case(32'h5fda3f91, 32'hdede1089);
	test_case(32'hdf6698f3, 32'hdde6dd74);
	test_case(32'hdfe10f48, 32'hdfe6d885);
	test_case(32'hdeda0f66, 32'hdfc0f9ba);
	test_case(32'hdff3ebd7, 32'hdfc54314);
	test_case(32'hdfe88fc4, 32'h5efbb7f5);
	test_case(32'hdecb8752, 32'h5ef421ed);
	test_case(32'hdfddfdaa, 32'hdf7efa24);
	test_case(32'hdecda7c9, 32'hdfe08b8d);
	test_case(32'hdec403b6, 32'hde419bc0);
	test_case(32'h5dc1238a, 32'hdff28b22);
	test_case(32'h5fc47142, 32'hde48bc66);
	test_case(32'hddf42744, 32'h5fe551bf);
	test_case(32'h5f545a5b, 32'h5fc82d94);
	test_case(32'h5f78f7ba, 32'hdfe5c1c0);
	test_case(32'h5f497a57, 32'h5fc81ad1);
	test_case(32'hdf700a32, 32'hdff3953c);
	test_case(32'h5fe5f732, 32'h5fe5e944);
	test_case(32'h5ef2efff, 32'h5f785c8c);
	test_case(32'hdd50bcdc, 32'hdfd4a7b3);
	test_case(32'h5f572a01, 32'hdecb44dd);
	test_case(32'h5fd864be, 32'h5f6d447d);
	test_case(32'hdff2ecc9, 32'h5fce0a24);
	test_case(32'hdfdfc0ed, 32'hdfdc9721);
	test_case(32'h5f606839, 32'hdffbd89e);
	test_case(32'hdffbf453, 32'h5fdf6d58);
	test_case(32'hdff8756e, 32'h5fe49ad2);
	test_case(32'hdec44489, 32'h5fe1ebfd);
	test_case(32'h5ec82ba5, 32'h5eefd9f6);
	test_case(32'h5ff8e9ea, 32'h5e4aa614);
	test_case(32'h5f6fe978, 32'hdfebaa84);
	test_case(32'hdeff12e9, 32'h5fe8f7f7);
	test_case(32'h5ff8809a, 32'hdfd14966);
	test_case(32'h5fc12669, 32'hdfc1ac52);
	test_case(32'h5f712ede, 32'h5fda6c17);
	test_case(32'h5f581f9f, 32'h5fcc01f7);
	test_case(32'h5fe5dcba, 32'h5ed912e4);
	test_case(32'h5fdfbebc, 32'hdff5aab3);
	test_case(32'hdf659e94, 32'hdfe93455);
	test_case(32'hdfd02f11, 32'h5ff81dfd);
	test_case(32'hdffddcc9, 32'h5f6cd9ac);
	test_case(32'h5d5efbfa, 32'h5ff9aa7c);
	test_case(32'hdf4d153f, 32'hdfcbf12f);
	test_case(32'h5f527cde, 32'h5e6c6a3f);
	test_case(32'hdfea1678, 32'h5ff51086);
	test_case(32'h5fcbb459, 32'hdfc9866b);
	test_case(32'hdf6deb5b, 32'hdf566fa9);
	test_case(32'h5ffc40c9, 32'h5fd682a1);
	test_case(32'h5fd264e1, 32'h5f67ff97);
	test_case(32'h5fded744, 32'hdfe74ce8);
	test_case(32'h5fe10afc, 32'hdfde46ce);
	test_case(32'hdd423af1, 32'hdf5035d4);
	test_case(32'hdfc3c5b9, 32'hdfc40db6);
	test_case(32'hde68a04f, 32'h5f7d5697);
	test_case(32'h5fc65bd1, 32'hdf445453);
	test_case(32'hdec197ec, 32'h5f5d6e30);
	test_case(32'h5ff3c639, 32'hdfc0f99c);
	test_case(32'h5e4f3cac, 32'hdfce75c2);
	test_case(32'hdff891be, 32'h5ff46e93);
	test_case(32'hded34920, 32'hdc5c22b1);
	test_case(32'hdfc4ce20, 32'h5f7dfb99);
	test_case(32'h5ff04368, 32'h5ff232d2);
	test_case(32'hdff1df2e, 32'hdecbe7b5);
	test_case(32'h5f7259d6, 32'h5fe4345a);
	test_case(32'hdfe0d2d0, 32'h5fdc5044);
	test_case(32'h5e7d7fcd, 32'hdff82bfd);
	test_case(32'hdffdc9af, 32'hdfe8136a);
	test_case(32'h5fc9d05f, 32'hdf709873);
	test_case(32'hdee6a452, 32'hdfde5915);
	test_case(32'hdf7b4dba, 32'h5f5dfa73);
	test_case(32'h5fe33b61, 32'h5f5847a3);
	test_case(32'h5ffd5184, 32'hdff562c4);
	test_case(32'h5f4f4737, 32'hdf628190);
	test_case(32'h5fff80b2, 32'h5f49fec8);
	test_case(32'h5f7dee02, 32'hdedc210b);
	test_case(32'h5fd30b7f, 32'h5df5938c);
	test_case(32'hdfc62cbd, 32'h5ff9c5fb);
	test_case(32'h5f7a8fc8, 32'hdfc109b5);
	test_case(32'h5dcfea27, 32'h5edcb017);
	test_case(32'h5fd86b88, 32'hdf47048f);
	test_case(32'h5ee3fddd, 32'h5fedb1b6);
	test_case(32'h5fed4b2f, 32'h5fca98f0);
	test_case(32'hdf414905, 32'hdfe27afc);
	test_case(32'h5f70e7fa, 32'h5fdfaff7);
	test_case(32'h5fc9e131, 32'h5fef442b);
	test_case(32'hded493f5, 32'h5ff97c79);
	test_case(32'hdfc34c42, 32'hddfb7a30);
	test_case(32'h5f61400e, 32'h5ff6762e);
	test_case(32'h5ffbb690, 32'hdfc65a06);
	test_case(32'h5fc33ae4, 32'h5fe615e6);
	test_case(32'h5f6edf9d, 32'h5e61c6c2);
	test_case(32'h5f4f5025, 32'h5ff72013);
	test_case(32'h5fee15ee, 32'h5fd8cf64);
	test_case(32'hdf721388, 32'h5f4e23c8);
	test_case(32'hde4f3980, 32'h5fcd6041);
	test_case(32'h5fe155ec, 32'h5fd24528);
	test_case(32'h5f66596a, 32'h5dd61051);
	test_case(32'hdf4ba72c, 32'hdfd4f39a);
	test_case(32'hdffd5ec1, 32'h5fc8f530);
	test_case(32'hdf5985d4, 32'h5fc7da2c);
	test_case(32'h5fecea25, 32'h5fcbd3b5);
	test_case(32'h5ffe053a, 32'h5d6446f0);
	test_case(32'hdedec9c5, 32'hdf63abbd);
	test_case(32'h5fdd80cb, 32'hdff87b12);
	test_case(32'hdfe25008, 32'h5ffee9b4);
	test_case(32'hde43da9c, 32'hdfd16e0d);
	test_case(32'h5fd752ed, 32'h5fd96c6b);
	test_case(32'h5f7faa05, 32'hded6007e);
	test_case(32'hdfd4adb0, 32'h5fccb89a);
	test_case(32'hdf68a5c8, 32'hdfcd8c33);
	test_case(32'h5f62f113, 32'h5eda15e0);
	test_case(32'h5fda07be, 32'hdfe08ebc);
	test_case(32'hdfececb0, 32'hdf5e9cf5);
	test_case(32'h5f49f78b, 32'hdf7d51e5);
	test_case(32'hde745573, 32'h5fcce4d4);
	test_case(32'h5fcd659d, 32'h5fcda90f);
	test_case(32'h5f755d64, 32'hdfe4b4fa);
	test_case(32'h5fc6a17d, 32'hdf5b6d1b);
	test_case(32'hdf415da8, 32'h5fc00a1d);
	test_case(32'h5f7193ca, 32'hdfd2e6b1);
	test_case(32'h5fffd1fa, 32'h5ffed6b3);
	test_case(32'hdfd177fa, 32'hde519aad);
	test_case(32'h5f441ad3, 32'h5ed30cae);
	test_case(32'h5ffe6119, 32'hdee5f231);
	test_case(32'h5ff2a0ec, 32'hdff6e2c7);
	test_case(32'hdfea2c22, 32'h5fdff051);
	test_case(32'hdffb37c2, 32'hdffd5daa);
	test_case(32'h5fcb51a9, 32'h5f724b5d);
	test_case(32'h5ef4956e, 32'h5fc3ede6);
	test_case(32'hdedb77cb, 32'hdef93b5f);
	test_case(32'h5e7f275d, 32'h5f63056b);
	test_case(32'h5ff3d872, 32'h5efce7bf);
	test_case(32'hdfd18bc3, 32'h5fc89333);
	test_case(32'hdef217d9, 32'h5fe8f327);
	test_case(32'h5f5a2620, 32'h5e7113be);
	test_case(32'h5fec613d, 32'hdee500dc);
	test_case(32'hdf408d7e, 32'h5fea0814);
	test_case(32'h5f7588e9, 32'hdfe0947e);
	test_case(32'h5feac821, 32'hdf7e5579);
	test_case(32'hddf71c7f, 32'hdf7ccfcd);
	test_case(32'h5ece2d13, 32'hdfe33caf);
	test_case(32'h5fda0c3c, 32'h5eca913b);
	test_case(32'hddcc791a, 32'hdf757af0);
	test_case(32'hde5af9b7, 32'h5e779e85);
	test_case(32'hdfe1182c, 32'hdfe10ad6);
	test_case(32'hdfee5b2d, 32'hdff9e0d5);
	test_case(32'h5ffa010f, 32'h5ee5accb);
	test_case(32'hdfd5c7be, 32'h5fd41ace);
	test_case(32'h5fe0c2c7, 32'hdfeb8cb6);
	test_case(32'h5f454ab7, 32'hdf50f1de);
	test_case(32'h5fdc3319, 32'h5fed382d);
	test_case(32'hdf4faca3, 32'hdf4ccd12);
	test_case(32'h5dce95a7, 32'h5ff45278);
	test_case(32'hdf6cb68d, 32'hdfc8caa1);
	test_case(32'hdedd5732, 32'h5f792ef7);
	test_case(32'h5f4788e1, 32'hdf6ffdef);
	test_case(32'hdb5000a1, 32'h5fc8f2ab);
	test_case(32'h5f607a8f, 32'hdfcda394);
	test_case(32'h5dfc10e3, 32'h5f46de0e);
	test_case(32'h5ed19c5c, 32'hdffe401b);
	test_case(32'hddd41aef, 32'hdfd943f9);
	test_case(32'hdf5e3110, 32'hdf75d600);
	test_case(32'h5f59eb19, 32'h5fea15cc);
	test_case(32'hdff7e23a, 32'hdfe3f408);
	test_case(32'h5ecc42cd, 32'hdfe82d17);
	test_case(32'hdfcaf909, 32'h5d50a769);
	test_case(32'h5f713e17, 32'hdcf4eb5d);
	test_case(32'hdfd8a244, 32'h5ed1f796);
	test_case(32'h5fd82946, 32'h5dcc7d00);
	test_case(32'h5fff9127, 32'h5feb61a8);
	test_case(32'hdfcd465b, 32'h5f4bac06);
	test_case(32'h5eefa88f, 32'hdfc7e74b);
	test_case(32'hded63f89, 32'hdef671be);
	test_case(32'h5fcf1cb5, 32'hdf5951c1);
	test_case(32'h5ffcc636, 32'hde78c691);
	test_case(32'hdf700710, 32'h5f4bc9a6);
	test_case(32'hdfe6b07b, 32'hdfe665a2);
	test_case(32'hdf60f06e, 32'hdf6e304c);
	test_case(32'h5f757f31, 32'hdfed37f2);
	test_case(32'h5e47abe2, 32'h5f4f2f3d);
	test_case(32'hdffebd2d, 32'h5fcadbd8);
	test_case(32'hdf42073d, 32'h5fe440b5);
	test_case(32'h5ff39df7, 32'hdfc4ab79);
	test_case(32'hdfc1831f, 32'hdee00398);
	test_case(32'h5ed3f004, 32'h5fc2fa80);
	test_case(32'hdfee40eb, 32'hdfefe92f);
	test_case(32'hdf7fa578, 32'hdf6b878f);
	test_case(32'hdfd45870, 32'h5f6eeb71);
	test_case(32'h5ee0e755, 32'h5ee57bb1);
	test_case(32'hdfc53c35, 32'h5ff9e8ed);
	test_case(32'h5f4d4998, 32'h5ee3c93f);
	test_case(32'hdcf527d9, 32'hdeefd828);
	test_case(32'hdfdd90d0, 32'hddce5619);
	test_case(32'hde6d27c1, 32'h5f77e13d);
	test_case(32'h5eedfaaf, 32'hdb56c817);
	test_case(32'hdeec7b4c, 32'hdfecc542);
	test_case(32'hdf4177e1, 32'hdfccb1b8);
	test_case(32'h5f5bde7c, 32'hdfdd01cd);
	test_case(32'h5fcdf1b7, 32'h5ecafc0a);
	test_case(32'h5f516eb2, 32'hde4b356d);
	test_case(32'h5ffa4645, 32'h5fe05ad6);
	test_case(32'hdefb63fd, 32'h5ec5525f);
	test_case(32'h5f406514, 32'hdec5dcd1);
	test_case(32'hdfe0b95c, 32'hdd63dc55);
	test_case(32'hdfecc3d7, 32'h5fc23acb);
	test_case(32'hdfeeb22c, 32'h5fedcef6);
	test_case(32'h5e42a8d9, 32'hdfeaaea5);
	test_case(32'hde6d793b, 32'hde71f43f);
	test_case(32'h5ffc4f96, 32'h5fe2878e);
	test_case(32'hde42e749, 32'hdfd59294);
	test_case(32'hdfdd2f04, 32'h5efae287);
	test_case(32'hded5df45, 32'hdef8730d);
	test_case(32'h5ec0210e, 32'h5f72f785);
	test_case(32'hdfd8a972, 32'hdffdaf4b);
	test_case(32'hdfce19a2, 32'hdff53603);
	test_case(32'hdec89014, 32'hde581d65);
	test_case(32'hdfcf8c8c, 32'h5f469fb0);
	test_case(32'hde6f9025, 32'hdf5a6a8c);
	test_case(32'h5e4f61dc, 32'h5fe5d8d1);
	test_case(32'hde63eb78, 32'h5fe7359a);
	test_case(32'h5c59a210, 32'h5fc3d7b9);
	test_case(32'hdff44379, 32'hde5fbeac);
	test_case(32'hded3c896, 32'hdf7966e7);
	test_case(32'hded3d6d0, 32'h5e5194c8);
	test_case(32'hdf6ad522, 32'hdfc72516);
	test_case(32'h5f54ff01, 32'hdf565013);
	test_case(32'h5eda3451, 32'hded01ae8);
	test_case(32'h5ffbce01, 32'hdf5182c9);
	test_case(32'h5fcd7097, 32'h5f79850f);
	test_case(32'hdefa24c2, 32'hdfc358dd);

    $finish;
end

task test_case(
    input [31:0] a_in,
    input [31:0] b_in
); begin
    @(negedge clk) begin
        a = a_in;
        b = b_in;
    end
    @(posedge clk) begin
        $display("%h,%h,%h", a_in, b_in, out);
    end
end
endtask

endmodule
