`timescale 1ps/1ps

`include "fadd.v"

module fadd_tb;

reg [31:0] a, b;
wire [31:0] out;

reg clk = 1'b1;

fadd uut(a, b, out);

always clk = #5 ~clk;

initial begin

	$dumpfile("fadd_out.vcd");
	$dumpvars(0, fadd_tb);
	test_case(32'hE0461BEC, 32'h5F0D7B6D);
	test_case(32'h5EA7FAD1, 32'hDF4C617E);
	test_case(32'hDFB6B9D2, 32'h5FBFBD16);
	test_case(32'hDF3B8DB3, 32'hDEB14EDE);
	test_case(32'hDFE6DD15, 32'hDECEF42A);
	test_case(32'h5F1323DA, 32'hDF745CFE);
	test_case(32'h5F775DF7, 32'hDEE5E075);
	test_case(32'h6070CC71, 32'h605ECB01);
	test_case(32'hDF3F607F, 32'h602A66C4);
	test_case(32'hDF791A4B, 32'h6011D200);
	test_case(32'h606FE34B, 32'hDF8EA64B);
	test_case(32'hE03E4C05, 32'hDFC97D63);
	test_case(32'hE01F876F, 32'hDEF9D073);
	test_case(32'h60657371, 32'h602F141B);
	test_case(32'hE02AF1BA, 32'h5F76D567);
	test_case(32'h5F44B445, 32'hDEE7AAB2);
	test_case(32'hDF9E496A, 32'h5F16369B);
	test_case(32'hE077EA08, 32'hE03D02FA);
	test_case(32'hDFDE3FAF, 32'h5FC9C1B4);
	test_case(32'h6006EE49, 32'hDE6D8272);
	test_case(32'h604876AF, 32'hE06B52DB);
	test_case(32'h606F8283, 32'hDEB28799);
	test_case(32'hDEF0F93A, 32'hE043234F);
	test_case(32'hE06B8192, 32'h605ECFA3);
	test_case(32'h60732094, 32'hDEC33C8A);
	test_case(32'h605E048C, 32'h604033BC);
	test_case(32'h605E6FEB, 32'hDF49BEB1);
	test_case(32'h6020BA34, 32'h5D72EDD6);
	test_case(32'hE01E6A87, 32'hE00CED3A);
	test_case(32'h5E872E66, 32'hE025AC07);
	test_case(32'h5F37FC7B, 32'h5FB2206F);
	test_case(32'h600CF810, 32'h60772CCD);
	test_case(32'h604C8E5E, 32'hE0506BE8);
	test_case(32'h5F8DF615, 32'h605DACA7);
	test_case(32'hDF23B1B0, 32'h5C0E3A07);
	test_case(32'hE07AD888, 32'h60284B1F);
	test_case(32'hDFDD1C93, 32'hDF19C71E);
	test_case(32'h604845A5, 32'h6007C5DA);
	test_case(32'hE05AFB4D, 32'hE019C935);
	test_case(32'h60631765, 32'hDF25DAAB);
	test_case(32'h5F9940D1, 32'hE0611B6B);
	test_case(32'h5EC4C5AC, 32'h5FF67562);
	test_case(32'h606E6AB3, 32'hE01A21F5);
	test_case(32'hDEA0B4B9, 32'h5F2B9498);
	test_case(32'h601A74F2, 32'hDF150AA6);
	test_case(32'h601C95F6, 32'h5DE7ECCE);
	test_case(32'h5F8BDB3F, 32'h6059386D);
	test_case(32'h5FF4630C, 32'hDF82C685);
	test_case(32'hE0348842, 32'hDDEDD443);
	test_case(32'h60741E90, 32'hE04BE8A2);
	test_case(32'hDFB22B2F, 32'hE07ADE59);
	test_case(32'hDF81021F, 32'h5FC7162F);
	test_case(32'h602DFE87, 32'h601720FE);
	test_case(32'h605E38DB, 32'h5FF9D813);
	test_case(32'hE0701FAE, 32'h5F09DED3);
	test_case(32'hE05DA747, 32'h606F4163);
	test_case(32'hDDE87913, 32'h600885CB);
	test_case(32'h603FE623, 32'h5EEDFA20);
	test_case(32'h60286462, 32'hE026385A);
	test_case(32'hDF10162E, 32'h605FCBF9);
	test_case(32'h5E92FE04, 32'h5EC6CA52);
	test_case(32'hE00102E2, 32'hE0452A4E);
	test_case(32'h605E247F, 32'h603350F6);
	test_case(32'hE032511A, 32'h5F61F887);
	test_case(32'hDE4F94EB, 32'h60339A38);
	test_case(32'h60118EB2, 32'hDF2E5850);
	test_case(32'hDFCB1CD3, 32'hE02B51F7);
	test_case(32'h607FF479, 32'h601913DF);
	test_case(32'h5E0945FA, 32'h601DD578);
	test_case(32'h5F610D53, 32'h5D1465DF);
	test_case(32'h5EBDCD1E, 32'h5FB4EB4A);
	test_case(32'hE0515F87, 32'h5FE0AE4D);
	test_case(32'h606CA8F7, 32'h607E8B3D);
	test_case(32'h5F5C0F7C, 32'hDFEE2F30);
	test_case(32'h5F9D963C, 32'h6058DA8A);
	test_case(32'hE02A3366, 32'h5FFA9C89);
	test_case(32'hDDBB3F01, 32'hDEC57393);
	test_case(32'h5FE285E7, 32'hDFA82062);
	test_case(32'hDE953B83, 32'h5FDB9E78);
	test_case(32'hE058CC79, 32'hE02F59B5);
	test_case(32'h60401CB9, 32'h5F998807);
	test_case(32'hE0282DC4, 32'h6077DBC0);
	test_case(32'hE00F3FD5, 32'h604F3A87);
	test_case(32'hE03669F8, 32'hDF7BF259);
	test_case(32'hDFE5BBDF, 32'h6036F49B);
	test_case(32'hE04F2A1F, 32'h60162744);
	test_case(32'hDFA325F7, 32'h5F891B6E);
	test_case(32'h60648B63, 32'h5EFFEC46);
	test_case(32'h606D806A, 32'hE03142F6);
	test_case(32'h5EBA897E, 32'hDEE221F4);
	test_case(32'h60179BBE, 32'h5F7D1F00);
	test_case(32'h5F770F43, 32'h5FA67529);
	test_case(32'h601552A3, 32'hE073D2B9);
	test_case(32'hDFF70800, 32'hDFBBB0CC);
	test_case(32'hDFD1CCDC, 32'h60446412);
	test_case(32'hDFE157FF, 32'hE0647834);
	test_case(32'hE01134F2, 32'h60038C36);
	test_case(32'hE0116D95, 32'hDF592A1D);
	test_case(32'hE015D08A, 32'hDE662F77);
	test_case(32'hDFF3C91C, 32'h6042B06A);
	test_case(32'hE033AF96, 32'h5FEE1FEE);
	test_case(32'hDF7D9ADD, 32'hDFC92908);
	test_case(32'hE00C1232, 32'hE06E5289);
	test_case(32'h5FC803F1, 32'h5FFF5228);
	test_case(32'hE005A617, 32'h5F00AD37);
	test_case(32'h606E3208, 32'h5FD05390);
	test_case(32'h5C665C3E, 32'h60580735);
	test_case(32'h5E8A54FF, 32'hDF003895);
	test_case(32'h5EB82DED, 32'h6023FC5F);
	test_case(32'hE03FFAEA, 32'hE05CF5B6);
	test_case(32'h603C6423, 32'hDEF6C44A);
	test_case(32'hDE17C068, 32'hDE6E4E1C);
	test_case(32'h6023DE8C, 32'h600137AE);
	test_case(32'h602482A1, 32'h6021ACA3);
	test_case(32'h6079F464, 32'hDEDB2B69);
	test_case(32'hDE89E759, 32'h5E53BE97);
	test_case(32'hDF95ED1E, 32'h5FACCADD);
	test_case(32'hDFDC1E66, 32'h5F2E4271);
	test_case(32'hE013B538, 32'hDED8EA2F);
	test_case(32'hE06FC224, 32'h5FBAF60C);
	test_case(32'hDFA21E99, 32'hE00AA468);
	test_case(32'h5F3A785B, 32'h60597224);
	test_case(32'h60297A14, 32'h5FF176C4);
	test_case(32'h5F85E345, 32'hE00C201A);
	test_case(32'hE0027998, 32'h5FF008D3);
	test_case(32'h607889F1, 32'h5D5C58A0);
	test_case(32'hE013F3B9, 32'hDF0248B4);
	test_case(32'hE0038A1C, 32'hE01A9351);
	test_case(32'hDF438078, 32'hDFF665F4);
	test_case(32'h5FAD262F, 32'h603BC12C);
	test_case(32'h5F9C29B8, 32'hDEBFE300);
	test_case(32'hDF2E0992, 32'h6031BB78);
	test_case(32'h5F0554C2, 32'h60028C54);
	test_case(32'h5FE18BB4, 32'hE026B3FA);
	test_case(32'h607A19F8, 32'hE045FB19);
	test_case(32'hE03CF8F4, 32'h6065BD3D);
	test_case(32'h6071F70C, 32'hDFE7C4D7);
	test_case(32'h5F212659, 32'hE0100E34);
	test_case(32'hDF9FC73E, 32'h5F347238);
	test_case(32'hDF6FE81C, 32'h5FC801E5);
	test_case(32'h5EE447D1, 32'h6009CB7F);
	test_case(32'h6054446A, 32'hE054605E);
	test_case(32'hDF9E184C, 32'hE0549AD1);
	test_case(32'h6032D718, 32'h60138C97);
	test_case(32'hE07B53EC, 32'hE064376C);
	test_case(32'hDF2284AB, 32'h5FDB2C50);
	test_case(32'hE05E2BD4, 32'hE07A0E1D);
	test_case(32'hDFFF815F, 32'hE00F2FF1);
	test_case(32'hE012B67D, 32'hDFE36C33);
	test_case(32'h5EE5E6D5, 32'h601AE90C);
	test_case(32'hDFAF496C, 32'h5EF898E8);
	test_case(32'hE07F8032, 32'h605BB99B);
	test_case(32'h5E878EA9, 32'h5FD0E46C);
	test_case(32'hDFCF30BA, 32'h6058963A);
	test_case(32'h5FC625FC, 32'h600796AC);
	test_case(32'h6029D8FA, 32'h6046140A);
	test_case(32'h6066DD61, 32'h5EA56EA7);
	test_case(32'hDFCC0A66, 32'hE032D0DC);
	test_case(32'hE005CDF0, 32'h5FEABE87);
	test_case(32'h5EDE15BA, 32'hDE92AC30);
	test_case(32'hDF8BB807, 32'h6060CD52);
	test_case(32'h5F9DF90F, 32'hE07898C8);
	test_case(32'hDF58661C, 32'hDF1940A8);
	test_case(32'h5F9F816E, 32'h5FB320BE);
	test_case(32'hDF19469E, 32'hDFF0A581);
	test_case(32'h5F671974, 32'hE04DE18A);
	test_case(32'h60380B83, 32'h6021889F);
	test_case(32'h5FE9D1F6, 32'h5F766A30);
	test_case(32'h606AAA99, 32'h5F293ED7);
	test_case(32'h5FF2BAE6, 32'hDFB52325);
	test_case(32'hDF9264F6, 32'h607DC4C7);
	test_case(32'h6075CAC7, 32'hE0625ED6);
	test_case(32'hDEEA78B1, 32'h60130683);
	test_case(32'h6015E392, 32'h5FE7636B);
	test_case(32'h5F4BE6B1, 32'h5FF02507);
	test_case(32'h601D9DD0, 32'h6056D4F4);
	test_case(32'hE0370B81, 32'h607CE355);
	test_case(32'h5F7C5ADE, 32'hE02A5AFE);
	test_case(32'h5CB5EF31, 32'h5F496CFD);
	test_case(32'h6009C60B, 32'hE01426BC);
	test_case(32'h5F0CE386, 32'hE03036DD);
	test_case(32'hDFB04325, 32'hE07DA5A4);
	test_case(32'hDF353390, 32'hDFF30B0D);
	test_case(32'h5EA60D30, 32'hE07C2C84);
	test_case(32'hDFEE16F9, 32'h5FFC9C34);
	test_case(32'h60656587, 32'hE052A885);
	test_case(32'hDF3ABF71, 32'hDFECF04F);
	test_case(32'hE01503B7, 32'hDF9CFCA9);
	test_case(32'hE027B115, 32'hDFC0E0A2);
	test_case(32'hE00BCEF0, 32'hDFCC180B);
	test_case(32'h5F5DD2E2, 32'h5ECE5E70);
	test_case(32'h601AB2BC, 32'hE049B60B);
	test_case(32'hDFA011D6, 32'hDFD35435);
	test_case(32'h600CD4D5, 32'hDFEC6E04);
	test_case(32'h6035EC4C, 32'hE06B8A1C);
	test_case(32'h60710DCA, 32'h604EEDDF);
	test_case(32'h5FFA2EAD, 32'h5D8CB1B5);
	test_case(32'hE03275EF, 32'h5F29F7B0);
	test_case(32'h604ACB9E, 32'hE059702D);
	test_case(32'hDF2A8B30, 32'h602F517A);
	test_case(32'h603E20D9, 32'h6023B1A3);
	test_case(32'h605856AB, 32'hDD43DF95);
	test_case(32'h5EE91BBA, 32'h601C7C5E);
	test_case(32'hDF9CCF0A, 32'h605CDCB0);
	test_case(32'hDFC698B7, 32'h5FB97A3E);
	test_case(32'hE0481283, 32'hE0422336);
	test_case(32'h5E0E0AC5, 32'hE01CF1F6);
	test_case(32'h5F372339, 32'h5FBCED17);
	test_case(32'h60191054, 32'h607C1E3C);
	test_case(32'h5F450A81, 32'hE003DE95);
	test_case(32'hE058E675, 32'hE03F3901);
	test_case(32'h5EDF5834, 32'h5AE07BD6);
	test_case(32'hE032FFA4, 32'hE07504B1);
	test_case(32'h5FD9AA50, 32'hE036ABF5);
	test_case(32'h5ED7AA24, 32'h60756A48);
	test_case(32'hE041232F, 32'h5E8405B2);
	test_case(32'hDEAE1388, 32'h5EEC7621);
	test_case(32'hDF3713F5, 32'h607E245D);
	test_case(32'hDF82DE9D, 32'hDEC57C8F);
	test_case(32'hE06835C9, 32'h5F63E94C);
	test_case(32'h5F8B1A94, 32'h5F93A1BB);
	test_case(32'h5F907897, 32'h5F4FAB53);
	test_case(32'hDF8DB928, 32'h5F832FBE);
	test_case(32'h60234770, 32'h606683A2);
	test_case(32'hDFA78BD6, 32'h60325764);
	test_case(32'h5EB6409A, 32'h6007B7DE);
	test_case(32'hDFB3E3BE, 32'h5F74098A);
	test_case(32'h5F26088B, 32'h6015434F);
	test_case(32'hE0051CBB, 32'h6006F57A);
	test_case(32'h5F0C9408, 32'hE07604FE);
	test_case(32'hDFD4717E, 32'hDE14703A);
	test_case(32'hE02CAB96, 32'hDF07B36F);
	test_case(32'hDFFD34DE, 32'h60558D3F);
	test_case(32'h5FEE9DA2, 32'h60643F35);
	test_case(32'h601D40B2, 32'h5FC5D5DA);
	test_case(32'hDFB58F64, 32'hDFE246DB);
	test_case(32'hE064F068, 32'h60656B62);
	test_case(32'hDFD2FBA8, 32'hE0330F8F);
	test_case(32'h604D860D, 32'hE0165923);
	test_case(32'hE05C86D6, 32'hE0761CA7);
	test_case(32'hE018638E, 32'h60556AB0);
	test_case(32'h5E23C6AE, 32'hDEF83C02);
	test_case(32'hDFDD0493, 32'hE0485FEC);
	test_case(32'h602C2DF9, 32'h60745549);
	test_case(32'h6059A6E4, 32'hE06085C3);
	test_case(32'hDFA9CB79, 32'hDFE5391C);
	test_case(32'hDF2031E1, 32'hE05E6B45);
	test_case(32'h5E90BEFD, 32'hDF8F32DF);
	test_case(32'hE02A49E0, 32'hE00BBA6E);
	test_case(32'hE0761071, 32'h601AA1D3);
	test_case(32'hE03B144D, 32'h6012A706);
	test_case(32'h6029F826, 32'hE0010EA9);
	test_case(32'hDF3F3FCC, 32'hE0390EBB);
	test_case(32'h5F0D2C47, 32'hE0768A13);
	test_case(32'hDF8CF72E, 32'h60657BBD);
	test_case(32'h5FCB50CE, 32'h600CF1EE);
	test_case(32'hE02D3817, 32'hDE0D9251);
	test_case(32'h5EF8AFA8, 32'h5F645516);
	test_case(32'h5F147C10, 32'hDF8DC45E);
	test_case(32'h605C9A67, 32'hE006345E);
	test_case(32'hDE046551, 32'h600EED79);
	test_case(32'h5EFD68EB, 32'hDFDBE7B0);
	test_case(32'hE0115AE4, 32'h5FC71C1B);
	test_case(32'h5F5C9B1C, 32'hE051BABE);
	test_case(32'hE0646A3D, 32'hE0132DDC);
	test_case(32'hDDAD81DB, 32'hE058A49A);
	test_case(32'hE0324558, 32'hE05D206C);
	test_case(32'h5EA44D83, 32'h60422A55);
	test_case(32'hDFBD1F3E, 32'hDFCE7719);
	test_case(32'h6065CDA0, 32'h5DB57ACE);
	test_case(32'hDF897587, 32'h5F3E20E2);
	test_case(32'hE07BEBA3, 32'h5FEC7C9C);
	test_case(32'hE04757FA, 32'hE050FAB6);
	test_case(32'h5FCC634B, 32'hDFA85D6C);
	test_case(32'h5F70A21A, 32'hE0169753);
	test_case(32'hE016AA8C, 32'h5EB7A6FF);
	test_case(32'hE0756D47, 32'hE071EFC5);
	test_case(32'h606C5FCC, 32'hDFFB3997);
	test_case(32'h5F9E1A78, 32'h600432EF);
	test_case(32'h5B7ACC8F, 32'hE061C56B);
	test_case(32'h607E04E7, 32'hE0059749);
	test_case(32'hE06C7D54, 32'h602BEFA4);
	test_case(32'h5FB06C7C, 32'h5F87EFF3);
	test_case(32'h600F3873, 32'h604CFE25);
	test_case(32'h60467B78, 32'hE052F46C);
	test_case(32'h60732199, 32'h6074CDA7);
	test_case(32'hDF9DA87B, 32'h5F3BD05C);
	test_case(32'h5E20544A, 32'hDE473892);
	test_case(32'hDE74A8E3, 32'hE06036CF);
	test_case(32'h5F283716, 32'hE04A34C5);
	test_case(32'hE00F85B5, 32'hDFA54745);
	test_case(32'h5F26F0A4, 32'hDF793CFF);
	test_case(32'h60133EE4, 32'h5F8F3807);
	test_case(32'hDFE0EE89, 32'hDF826F6F);
	test_case(32'h5D7F9EF1, 32'h600AA139);
	test_case(32'h5ED3B1CA, 32'hDF4A2369);
	test_case(32'h5E80EF30, 32'hE00A1DB8);
	test_case(32'h607D8BF7, 32'h606865EF);
	test_case(32'h5F3D2078, 32'hDF3638FC);
	test_case(32'h60646A1A, 32'hDE03633A);
	test_case(32'hE00179CC, 32'hDF98D199);
	test_case(32'h6058DD0E, 32'h5FD7EFB0);
	test_case(32'h6016A1AE, 32'hE03DE409);
	test_case(32'hE07B7A13, 32'hDF528CD0);
	test_case(32'h5FD3676E, 32'hE03ED5D0);
	test_case(32'h605B4127, 32'hE03D1D49);
	test_case(32'h5D9055CF, 32'h6011B398);
	test_case(32'hE0203CEC, 32'hE05CF525);
	test_case(32'h5EBD6B5D, 32'h5FBA8524);
	test_case(32'hDE48C2DC, 32'h60321B98);
	test_case(32'h6034083B, 32'h6065F5CF);
	test_case(32'h5F9573EB, 32'hDF0F082B);
	test_case(32'h5F569211, 32'h6029EF81);
	test_case(32'hE05002AF, 32'h605AF5BE);
	test_case(32'hE00746B5, 32'hDEC9B58D);
	test_case(32'h5FAC07D8, 32'h5FFB7D1E);
	test_case(32'h5DB6301B, 32'h6059CE8D);
	test_case(32'hDFE27615, 32'h5FC61149);
	test_case(32'hE003BEE9, 32'hE00EF115);
	test_case(32'hE0133B53, 32'h601AFEC9);
	test_case(32'h5FCC1ACA, 32'h5FEFAA21);
	test_case(32'hE03EBF2C, 32'hDF4AB8D1);
	test_case(32'h5F99F634, 32'h605FEF55);
	test_case(32'h5ECB5778, 32'hE033CFE2);
	test_case(32'hDFCA6B82, 32'hDF189F95);
	test_case(32'hDE2993D0, 32'h5E4EC85C);
	test_case(32'hDFE41EFC, 32'h6042D84B);
	test_case(32'hDFE8A7AA, 32'h602E42B0);
	test_case(32'hE05E6520, 32'hDFBBBBD5);
	test_case(32'hE018ADE4, 32'hDFA7869E);
	test_case(32'h5F292DB4, 32'hDF1F71A2);
	test_case(32'h5FF3B430, 32'h5FD90ED3);
	test_case(32'h5F8F2BFF, 32'h605E74FD);
	test_case(32'hDFEC9D46, 32'hE077915C);
	test_case(32'hDFA4D2E4, 32'hDE96E6E1);
	test_case(32'hDF5C54E8, 32'h5FAF1C6B);
	test_case(32'h6007E5E6, 32'hE06E79F7);
	test_case(32'h604EB6C0, 32'h6030281B);
	test_case(32'h5D8B090D, 32'h60171E0E);
	test_case(32'hE059C684, 32'h602CB78D);
	test_case(32'hDFB4FDCB, 32'hDE878B12);
	test_case(32'h607537B3, 32'hDF74AFB9);
	test_case(32'hE0294345, 32'hDFC8E024);
	test_case(32'hE0241373, 32'h5FFD7361);
	test_case(32'hDDD295FB, 32'hE04C9D72);
	test_case(32'h606200C1, 32'h6055A7AD);
	test_case(32'hDECC4D3E, 32'h5F876706);
	test_case(32'h60027AD9, 32'h5FD754E9);
	test_case(32'hE07A75C9, 32'hDF8F1CDC);
	test_case(32'hE0713E22, 32'h6045F760);
	test_case(32'h604A1469, 32'hE0713EB5);
	test_case(32'h603C394D, 32'hE0328DB1);
	test_case(32'h60057B9F, 32'h607212CF);
	test_case(32'h603CF39B, 32'hE02BA4A9);
	test_case(32'h6031D434, 32'hDF4AC206);
	test_case(32'hE061E356, 32'hDF9828CF);
	test_case(32'hDFEE0F05, 32'hE069B395);
	test_case(32'hDFEDA340, 32'h5FE8B31F);
	test_case(32'h6032514B, 32'h602FE16B);
	test_case(32'h6053C133, 32'hE070D109);
	test_case(32'hDEF4B80D, 32'hE048C261);
	test_case(32'h5F63E8F5, 32'h604F03F4);
	test_case(32'h5FEC2C4B, 32'h60734DF4);
	test_case(32'h5F0DE6B0, 32'hE02F6C46);
	test_case(32'h606ADA0F, 32'hDF3462B0);
	test_case(32'h5FDDCE02, 32'hDFBFFFAA);
	test_case(32'hDFD04DD2, 32'hDFB8F823);
	test_case(32'hE070BECC, 32'hE07CF0BB);
	test_case(32'hE026AD6B, 32'hE03CD4E8);
	test_case(32'hE02F6788, 32'hDD28CF11);
	test_case(32'hDF805EEE, 32'hE00A1CC0);
	test_case(32'h6074FB10, 32'h5FFADBB6);
	test_case(32'hDF426108, 32'hDEEF006F);
	test_case(32'hDED0790B, 32'h60314A60);
	test_case(32'hE05D054B, 32'h602773A0);
	test_case(32'hE053C476, 32'h602A517A);
	test_case(32'h5E3CE99F, 32'hE04815E5);
	test_case(32'h5FA82FDC, 32'h602EF95D);
	test_case(32'hDFEF27F7, 32'hE020D939);
	test_case(32'h5FB1CCAE, 32'hE0443E59);
	test_case(32'h6009C017, 32'hE03740DA);
	test_case(32'h606EADAF, 32'h5F13DD41);
	test_case(32'h6052766E, 32'h60055489);
	test_case(32'hDF3B2E09, 32'h5FA9C4C8);
	test_case(32'h603358C9, 32'h601C60F4);
	test_case(32'h606F92D7, 32'h603F1B2B);
	test_case(32'h6012922C, 32'hDF928D27);
	test_case(32'hDFDE574A, 32'h60237C85);
	test_case(32'h6024021A, 32'h5ED47951);
	test_case(32'hE05FBD94, 32'hDFB307DE);
	test_case(32'hE043F3A1, 32'h5F1D3C0A);
	test_case(32'hE01EA465, 32'hDFDA453F);
	test_case(32'h5F9B139A, 32'hE006D982);
	test_case(32'h5FC74548, 32'hE0197967);
	test_case(32'hE05A1F63, 32'h601FA1E0);
	test_case(32'hE048C270, 32'h5FD69E44);
	test_case(32'h5F14E9CC, 32'h5F457241);
	test_case(32'h5FBDBAFD, 32'h5F8D4D78);
	test_case(32'h601A0898, 32'h601A0D45);
	test_case(32'hE0626169, 32'hDFBC9210);
	test_case(32'hE06A4347, 32'h605165B7);
	test_case(32'hE0059C4C, 32'h5F73C9D8);
	test_case(32'h601F1E02, 32'h605D639F);
	test_case(32'h60316440, 32'h5FD0AA48);
	test_case(32'hDFB94E80, 32'h5F9A7F8A);
	test_case(32'h601C184A, 32'hDF75D2E2);
	test_case(32'h5F95C930, 32'hE053B1A8);
	test_case(32'h5EF00E62, 32'h6049C18E);
	test_case(32'h5FE1804A, 32'h6041A093);
	test_case(32'hDF860475, 32'h605EEFBD);
	test_case(32'h602C78E5, 32'hDFEE214C);
	test_case(32'h60251078, 32'h604E223C);
	test_case(32'hDED4AB7C, 32'hDEC33672);
	test_case(32'hE0710DDC, 32'h60270000);
	test_case(32'hDF774E38, 32'hDFADEFEE);
	test_case(32'hE02C1DBD, 32'hE03490DD);
	test_case(32'hE0018A47, 32'h5E2B8B6C);
	test_case(32'h6015584A, 32'h603591B4);
	test_case(32'h5E9D701B, 32'h60724682);
	test_case(32'hE00E188D, 32'h5CCCB162);
	test_case(32'h5FEE6751, 32'hE059E382);
	test_case(32'hDF822110, 32'hE036A049);
	test_case(32'hDFEC61F1, 32'h5E2B2759);
	test_case(32'h5FA078EE, 32'h5E90343E);
	test_case(32'h5F24D242, 32'hDF650707);
	test_case(32'hE00603A0, 32'h604E7D0D);
	test_case(32'h5F4080F9, 32'h606A0475);
	test_case(32'h600B8EEC, 32'hE04F8059);
	test_case(32'h601342C6, 32'hE07B1DF9);
	test_case(32'hE025D826, 32'h5F20248F);
	test_case(32'h60387A1D, 32'hE05678F9);
	test_case(32'h606AFD64, 32'h5F3CDFFC);
	test_case(32'hE031A3FC, 32'h606ECF6A);
	test_case(32'h605E48D0, 32'hDE25C78A);
	test_case(32'h605F30F1, 32'h5DE46F4E);
	test_case(32'h5F34D55A, 32'h6055FC8E);
	test_case(32'h5FEABAB1, 32'hE0514C3C);
	test_case(32'hDEA6E023, 32'h5FD8A8FD);
	test_case(32'hDF99B709, 32'hE030916E);
	test_case(32'h60035D0F, 32'hDF2226B5);
	test_case(32'hE05AED1A, 32'hDFE6CD00);
	test_case(32'hE004C65F, 32'h5F583E8F);
	test_case(32'hDFB8C56C, 32'h5EEC9D40);
	test_case(32'hE06A68A5, 32'hDFC2AC11);
	test_case(32'hE0228ADD, 32'h6037677D);
	test_case(32'hE02BACC3, 32'h5EAC9C8F);
	test_case(32'h5ECBFFA1, 32'h5F277BC9);
	test_case(32'h6027109D, 32'h607B9127);
	test_case(32'h5EC6F96D, 32'h606063FC);
	test_case(32'hE013676B, 32'hDFAD0B8A);
	test_case(32'hDEE4E3C6, 32'hE030351E);
	test_case(32'hDF907747, 32'h5F930B87);
	test_case(32'hDD48B745, 32'hDDF8C02A);
	test_case(32'h5F02956C, 32'h6066DD31);
	test_case(32'h5F182223, 32'hDF0B4900);
	test_case(32'hDFA3CFF4, 32'hE03B70D8);
	test_case(32'h5F86E524, 32'hDE531495);
	test_case(32'h5FB3157E, 32'hE015F6B6);
	test_case(32'h5FCD0E43, 32'h5EE55D0F);
	test_case(32'hE032DAA8, 32'h601839CB);
	test_case(32'h60666043, 32'h603E946C);
	test_case(32'hE0647EB9, 32'hDF5898FB);
	test_case(32'h6017B30C, 32'hE045D15C);
	test_case(32'hDF4A8A8C, 32'hDFAFE35A);
	test_case(32'hE064201D, 32'h5F97AF77);
	test_case(32'hE05DE738, 32'h5EEBD51A);
	test_case(32'h600EE97A, 32'h603C363B);
	test_case(32'hDFD6A00D, 32'hE0424143);
	test_case(32'hE02F91E9, 32'h5E929FEC);
	test_case(32'hDFCBF97D, 32'h5F909C7D);
	test_case(32'h60214077, 32'h5E8210C1);
	test_case(32'h5FDF3E62, 32'h60194837);
	test_case(32'hE04CD011, 32'hE01FE78E);
	test_case(32'h6063A6F1, 32'h6033BC90);
	test_case(32'hDF14D832, 32'h6027F238);
	test_case(32'h5FE636DC, 32'hE015B6AA);
	test_case(32'h606C3C82, 32'h5FA71F30);
	test_case(32'hDFF096B0, 32'hDF9529DA);
	test_case(32'h5F8A222D, 32'h607121A3);
	test_case(32'h5FA1E191, 32'h5F64BF16);
	test_case(32'hE0387CFB, 32'h6037CF88);
	test_case(32'h601C6105, 32'hE017DF16);
	test_case(32'h5F83B7C6, 32'hDF83B051);
	test_case(32'hDFF0B1B0, 32'hDF78C362);
	test_case(32'h6002554E, 32'hDE2CB531);
	test_case(32'h5FB3B167, 32'h60744E0D);
	test_case(32'hE027A3BF, 32'hDFC552F8);
	test_case(32'hE0307BF5, 32'h605A3A4D);
	test_case(32'hDF64A524, 32'h6040ABCB);
	test_case(32'h5FBB165B, 32'hDED1EE6D);
	test_case(32'h5FD10348, 32'h60212C67);
	test_case(32'hE0488827, 32'hE0032D5F);
	test_case(32'h600F39CB, 32'hDF72FD6B);
	test_case(32'h60496547, 32'hDE46ECA0);
	test_case(32'h602C79C7, 32'h60548ADA);
	test_case(32'h5F9ECE43, 32'hE0091CD4);
	test_case(32'hE00BEDB7, 32'h604AE2EB);
	test_case(32'h5F942C2A, 32'h605EB566);
	test_case(32'hE007DCA0, 32'h603488CC);
	test_case(32'hDF8E668C, 32'h5F43BC4F);
	test_case(32'h5F160D17, 32'h607EADEA);
	test_case(32'hE058D873, 32'hDEE9E13A);
	test_case(32'hDDF75A80, 32'hE0634A31);
	test_case(32'h5EBA80C0, 32'hDF6A75F0);
	test_case(32'h607A36F5, 32'hDF8B059B);
	test_case(32'hDFE61F0D, 32'hDE594F95);
	test_case(32'h6016AAE0, 32'h5FDB059B);
	test_case(32'h606B2494, 32'hE0153332);
	test_case(32'h5D88257E, 32'h6024F2EB);
	test_case(32'h60655C5B, 32'h607E6FBC);
	test_case(32'h6000394A, 32'hDF52C490);
	test_case(32'h60027767, 32'h601859B7);
	test_case(32'hDF0CE8B9, 32'hE07D715A);
	test_case(32'h5F2126F8, 32'h5F2562A6);
	test_case(32'h5F0A50DB, 32'h604DC8CD);
	test_case(32'hDE6FE4F4, 32'hE0765B52);
	test_case(32'hDE2F04DF, 32'h5E7DFAEC);
	test_case(32'h60014683, 32'h5EFF6AE0);
	test_case(32'hE01B2EC5, 32'hE03D43FA);
	test_case(32'hDF1E902C, 32'h5FFD8D3B);
	test_case(32'h5FD0C420, 32'hE07800D7);
	test_case(32'hE01D4475, 32'h5D2F5B32);
	test_case(32'hDEEF80CA, 32'h5FD83FAD);
	test_case(32'h6027C701, 32'h607AFE7A);
	test_case(32'hE030D475, 32'h600139B0);
	test_case(32'h603A250B, 32'h604A3831);
	test_case(32'h5F8755FE, 32'hDFB912EF);
	test_case(32'h5FA66565, 32'hDF085554);
	test_case(32'h5F330F35, 32'h606B7261);
	test_case(32'hE06D18F4, 32'h5F0B57F5);
	test_case(32'hDEEF3D26, 32'h5FAEA5B2);
	test_case(32'hE074CEB8, 32'h5EACEB50);
	test_case(32'h601CB6A0, 32'hE003A38E);
	test_case(32'hE05F61F1, 32'hE030397F);
	test_case(32'hE01743ED, 32'h6015737D);
	test_case(32'h5E5AA089, 32'h5EFFAB7A);
	test_case(32'hDF9EC273, 32'hE06DDDD0);
	test_case(32'h600EBAFE, 32'hE011C1A3);
	test_case(32'h5E46CDD3, 32'hE0746F95);
	test_case(32'h5D0EFD84, 32'hDF67650B);
	test_case(32'h6005432C, 32'hDFC9805B);
	test_case(32'h5FD78755, 32'hDF526872);
	test_case(32'h6001D47F, 32'hE011D307);
	test_case(32'h6047BFDC, 32'h5FD5B0B5);
	test_case(32'h5FC9CA6F, 32'hE015F340);
	test_case(32'h6078FC9D, 32'hDFC90396);
	test_case(32'hE00E6B59, 32'hE02434E4);
	test_case(32'hE010B2F0, 32'hDF843C53);
	test_case(32'hE03C7B23, 32'h603B5645);
	test_case(32'hDF059A0F, 32'hDF2A6B93);
	test_case(32'h6056B213, 32'hDF5B0B6F);
	test_case(32'h5EA9E944, 32'h5F3E967C);
	test_case(32'h607A7165, 32'h6046DD92);
	test_case(32'h5FF8060D, 32'hE02240D2);
	test_case(32'h601FE28B, 32'hE0621920);
	test_case(32'h6055347A, 32'h60378637);
	test_case(32'h5CF69EB9, 32'h5E5ECB26);
	test_case(32'hDFCF2EBC, 32'h601C428D);
	test_case(32'h6010E3F6, 32'hDB04852D);
	test_case(32'h5FBB1250, 32'hE01B487E);
	test_case(32'h605DD0AE, 32'hDF82BEB5);
	test_case(32'h5F441FDF, 32'h6071ACE3);
	test_case(32'h5F12BA39, 32'hDD9B5D9A);
	test_case(32'h5F1A3C40, 32'hE02D596B);
	test_case(32'h5F9B75D3, 32'h606774DD);
	test_case(32'hDEDD48C8, 32'hE00A2140);
	test_case(32'h600C6D63, 32'h605B7974);
	test_case(32'hDFC1A5D8, 32'h6036DFFB);
	test_case(32'hE07C1D60, 32'hE008488C);
	test_case(32'hE07263A6, 32'h5F36EB1D);
	test_case(32'hE07612A2, 32'h6035B8B5);
	test_case(32'h5FBB85D3, 32'hE03F1EEE);
	test_case(32'h5FAF6FDA, 32'hDF5D4FCC);
	test_case(32'h5F8D1797, 32'h5FFAE113);
	test_case(32'h5FF7D4A2, 32'h5E906CB6);
	test_case(32'hE03CAC7F, 32'h6071E656);
	test_case(32'h5E7BCFF3, 32'h5DDEDEE5);
	test_case(32'hE00F59C2, 32'h603F3090);
	test_case(32'h6024D5C8, 32'hE00C0F4A);
	test_case(32'hDF98E673, 32'hDE1AE525);
	test_case(32'hDFCE9C37, 32'hDFCD41B5);
	test_case(32'h602E0E25, 32'hE029DE1C);
	test_case(32'h5FDAFFAC, 32'h60375005);
	test_case(32'hDF2BB4E6, 32'h5FEAC6BE);
	test_case(32'h600CA9F2, 32'hE012916C);
	test_case(32'hE01195C7, 32'hDF2C1A03);
	test_case(32'h607CC18B, 32'hDEE16C80);
	test_case(32'h607EAABD, 32'h5FC27B05);
	test_case(32'hE042F91E, 32'h601BE88B);
	test_case(32'h606096EC, 32'h604F0751);
	test_case(32'hDFACA728, 32'h5F9ED0E5);
	test_case(32'hE04417C0, 32'hE001312A);
	test_case(32'h60165909, 32'h6056F5F5);
	test_case(32'hE048D7B9, 32'hDEE8FB33);
	test_case(32'hE016B06E, 32'h606D98B1);
	test_case(32'h5F0D2619, 32'hE01ECD3C);
	test_case(32'hE041C2E8, 32'h6058A514);
	test_case(32'hDEAC245D, 32'h60342293);
	test_case(32'h5FAA71FA, 32'hE0184B6A);
	test_case(32'h6011EE84, 32'h5F94A8A6);
	test_case(32'h603D972F, 32'hE0604CB5);
	test_case(32'hDF6EDC3A, 32'h5F553567);
	test_case(32'hDE566671, 32'hDFDA5916);
	test_case(32'h5FAF1B9B, 32'h600740A2);
	test_case(32'hE06281FA, 32'h60522BAB);
	test_case(32'hE03B59E5, 32'h5F787DC1);
	test_case(32'hE02C1036, 32'h607B02E8);
	test_case(32'h60192933, 32'hE0217C8F);
	test_case(32'hE0205F67, 32'hDFB2CDD2);
	test_case(32'h5E7EEBE2, 32'h6079C711);
	test_case(32'hE058790A, 32'h5E66E2D5);
	test_case(32'hE01DCC3B, 32'hDF7230B6);
	test_case(32'h60729F2C, 32'hDECB19E2);
	test_case(32'h5FBAB3BB, 32'hE007CD84);
	test_case(32'h605883B7, 32'hDFE89476);
	test_case(32'h601F4024, 32'hDFCD9353);
	test_case(32'h606E6D91, 32'hDE449CEB);
	test_case(32'hDFB8D3F7, 32'h5FA376C6);
	test_case(32'h603FB194, 32'hDFFCDDE4);
	test_case(32'h5F59DFAD, 32'h601277B3);
	test_case(32'hE00876EC, 32'h604656CE);
	test_case(32'hDFCE1FD9, 32'hDFF8F747);
	test_case(32'hE01A3495, 32'h5E7BB201);
	test_case(32'h600EFE65, 32'h601D9D64);
	test_case(32'hDFE14FF0, 32'h5F3FEE78);
	test_case(32'h5FB3EEE7, 32'h5F71B3E1);
	test_case(32'h600D77B7, 32'hE00CF8D5);
	test_case(32'h5F753CD8, 32'hE05AB27C);
	test_case(32'h5F88CC98, 32'hE056CB78);
	test_case(32'h600EDA5D, 32'h5FA24B3E);
	test_case(32'h5F15EE1A, 32'h60338720);
	test_case(32'hDF146B93, 32'h5FBAA276);
	test_case(32'h606198A1, 32'h60516183);
	test_case(32'h5E5097F5, 32'h5EA9E6CD);
	test_case(32'hDF79A0DB, 32'hDFDB67A8);
	test_case(32'hE010BFCF, 32'hE05FB486);
	test_case(32'h60217F68, 32'hE07B831E);
	test_case(32'h6044C2F4, 32'hE00E7FD0);
	test_case(32'h602F4598, 32'hDFB3536A);
	test_case(32'hDFCAFE55, 32'hE024E440);
	test_case(32'hDF2FC38D, 32'h5F806E02);
	test_case(32'h5F849EB0, 32'h6003C385);
	test_case(32'h5EF544D1, 32'h601614FF);
	test_case(32'h5FB98009, 32'h604827FC);
	test_case(32'h5F9E3BF7, 32'hDFBEB4CE);
	test_case(32'hE003F27A, 32'hE06CD50F);
	test_case(32'hE0099EE0, 32'hDFEF9394);
	test_case(32'hE06377EB, 32'hDFCEC334);
	test_case(32'h5FBCF8C4, 32'hDF1C6A64);
	test_case(32'h6046CF75, 32'hDEBE457D);
	test_case(32'h5FCCAFD5, 32'h5F763847);
	test_case(32'h605A954E, 32'hDDB657A0);
	test_case(32'h5DE533BA, 32'hE066558A);
	test_case(32'h5F8208F4, 32'hE0426894);
	test_case(32'h606184E5, 32'hE061BF00);
	test_case(32'hE077F157, 32'hE05BC39C);
	test_case(32'h5E52386A, 32'h6054EE70);
	test_case(32'h5FF08239, 32'hE07DE48F);
	test_case(32'h606AEF82, 32'hDFF0514B);
	test_case(32'hE01D9563, 32'h5FFC3988);
	test_case(32'hDF008CD4, 32'h5F74A0B9);
	test_case(32'hE074C775, 32'hE0462C88);
	test_case(32'hDEC80098, 32'hDF746D8B);
	test_case(32'h6041A4CF, 32'hDFD91885);
	test_case(32'hE0070B42, 32'hE00BD477);
	test_case(32'hDFCA31BB, 32'h5E9B0684);
	test_case(32'h605005DC, 32'hDF94F77C);
	test_case(32'h5FB34653, 32'h5ED501DC);
	test_case(32'h5FA8D31B, 32'h6074FA70);
	test_case(32'hDEAFC6C5, 32'hDFFB02ED);
	test_case(32'hDF8B77A7, 32'hDF9EF53D);
	test_case(32'h5FC24E71, 32'hE05B8F54);
	test_case(32'h60334DC3, 32'hDF81D767);
	test_case(32'hDFDC381D, 32'h5F5DD65D);
	test_case(32'hE067BD94, 32'hE041F187);
	test_case(32'h5FE42465, 32'hDFBCF721);
	test_case(32'hE001290D, 32'h6023BCE3);
	test_case(32'h5FC895E9, 32'hDFEA2039);
	test_case(32'h6000A318, 32'h5F588D70);
	test_case(32'hE00A76A2, 32'hE0513ECF);
	test_case(32'h5F5E3C3E, 32'hDEFEB2F5);
	test_case(32'hE01EB57D, 32'hDFB127CC);
	test_case(32'hE028A7CE, 32'hDF9874F8);
	test_case(32'h607523A4, 32'hE060C846);
	test_case(32'h5F526758, 32'h6055F9D8);
	test_case(32'hDD9ECBFB, 32'hDF8214DA);
	test_case(32'h603D10A3, 32'hE0136134);
	test_case(32'hE04A1967, 32'hE07BFA6D);
	test_case(32'h5F1CD413, 32'hE0066082);
	test_case(32'hDF8BA13E, 32'h607681D5);
	test_case(32'hDF1D6748, 32'hDFBF00E4);
	test_case(32'h5F0437B8, 32'h60675473);
	test_case(32'h6011009B, 32'h5E710ED8);
	test_case(32'hDFC96978, 32'h60758592);
	test_case(32'hDF3BF9C4, 32'hE024FE2B);
	test_case(32'hE0052EB1, 32'hDF88DDE1);
	test_case(32'hDFC86616, 32'h605CB6AA);
	test_case(32'h5F207073, 32'h5F471B36);
	test_case(32'hDFBC392F, 32'hDE526CCD);
	test_case(32'h607FAD21, 32'hE01B068B);
	test_case(32'hDEFB6B07, 32'hDDE310F2);
	test_case(32'h5EFE5D35, 32'h602BE521);
	test_case(32'hE05CBBFE, 32'h5FA3BC44);
	test_case(32'h5FA06541, 32'hDFF9C9F6);
	test_case(32'hDF881EEF, 32'h5FBE8CB2);
	test_case(32'hDFDC135B, 32'hDFE58373);
	test_case(32'h603BF923, 32'h6017B4CC);
	test_case(32'hE038798C, 32'h6025C85D);
	test_case(32'h603DF939, 32'hDDCC7B8C);
	test_case(32'hE0400F96, 32'hE03A7150);
	test_case(32'h5FA445CB, 32'hDF9ECC40);
	test_case(32'h606F86A7, 32'hDF46CDFD);
	test_case(32'hDEC35DD0, 32'h5FF32EA3);
	test_case(32'hDFF8E9A9, 32'h5EF8F1A3);
	test_case(32'hDFB7A3C1, 32'h5F880934);
	test_case(32'h5FCC3A21, 32'h60758751);
	test_case(32'h6050ECD8, 32'hE05487D0);
	test_case(32'h5F9278A6, 32'hE007A664);
	test_case(32'hDF360A15, 32'hE01A8420);
	test_case(32'h5FC02907, 32'hDF8C477D);
	test_case(32'h607377C8, 32'hDF243137);
	test_case(32'h607E6FDF, 32'hDF1D555A);
	test_case(32'h5E240148, 32'hE06831B1);
	test_case(32'hE077F19C, 32'h606B33AF);
	test_case(32'h605272C0, 32'h607ED92C);
	test_case(32'h60109398, 32'h6022DD32);
	test_case(32'hDFE0D650, 32'hDF0C3B99);
	test_case(32'hDFCDD7BB, 32'hE06F4765);
	test_case(32'hDFD34068, 32'hDFE13D7C);
	test_case(32'hE0020467, 32'hDE941C48);
	test_case(32'hE01287E1, 32'h5FEA246A);
	test_case(32'hE060C6AA, 32'h60748E7E);
	test_case(32'h607FBF60, 32'hDF1D5E4D);
	test_case(32'h600BF6DA, 32'hE014C40E);
	test_case(32'hDEADB79B, 32'h5FF6B3AD);
	test_case(32'h5F868A00, 32'hE055A5B2);
	test_case(32'h60630329, 32'h603EA8FD);
	test_case(32'h602A9405, 32'h5F1409D7);
	test_case(32'hDFB0D308, 32'h60224B5F);
	test_case(32'hDF983F26, 32'h601E90B5);
	test_case(32'h5FD1E7E3, 32'hE07C25DC);
	test_case(32'hDEA5ADEC, 32'h6023ECC3);
	test_case(32'h60082698, 32'hE00E7618);
	test_case(32'hE0542BC9, 32'h5F5EB6DF);
	test_case(32'hE029C5FD, 32'hDFC1D8B0);
	test_case(32'h6055BC75, 32'hDED6C081);
	test_case(32'h5FA27280, 32'hDF35760E);
	test_case(32'hE06E3940, 32'hDEA00E90);
	test_case(32'hE0647EA7, 32'hE03ECA07);
	test_case(32'h5EF204A4, 32'hDE8437EC);
	test_case(32'hDF1D2C3C, 32'hE05773B0);
	test_case(32'h5F310524, 32'hDF0A701D);
	test_case(32'hE0010AD2, 32'h5F254B9E);
	test_case(32'h5FC46A43, 32'hE07E8424);
	test_case(32'hDFB7B493, 32'hDFD51402);
	test_case(32'h5C8AB041, 32'hE029F64F);
	test_case(32'h5FEDA063, 32'hDDB10DA2);
	test_case(32'h6054038B, 32'h60261718);
	test_case(32'h606EA44D, 32'hDE02CE13);
	test_case(32'hE02A73CB, 32'hE00E5B8A);
	test_case(32'hE0618D8A, 32'hDE9B7E32);
	test_case(32'h5F2FA653, 32'h5F1BEC23);
	test_case(32'hDE9A6030, 32'hE03F65F0);
	test_case(32'hDF9A3FBA, 32'h600FFFBB);
	test_case(32'hDFC987BD, 32'h6014D39D);
	test_case(32'hDF44FF23, 32'hE06A36A2);
	test_case(32'h605F167E, 32'hE0420AFF);
	test_case(32'hDF943595, 32'hDF740731);
	test_case(32'hE0583A86, 32'h5F72776D);
	test_case(32'h5F1F79D6, 32'hE018E948);
	test_case(32'h60347F23, 32'hDF3C2112);
	test_case(32'hDFCD31E6, 32'hDE4DBAE9);
	test_case(32'hE0421E91, 32'hE04DB10B);
	test_case(32'hDF341ECC, 32'hE001F374);
	test_case(32'hE067D7AE, 32'hE00A8628);
	test_case(32'hE0511F89, 32'h5F776FEB);
	test_case(32'hDF170EA4, 32'h5F6843DB);
	test_case(32'hE03BFB55, 32'hDFFDF449);
	test_case(32'hDF1B4F92, 32'hE041171A);
	test_case(32'hDF08076D, 32'hDE833781);
	test_case(32'h5E024714, 32'hE0651645);
	test_case(32'h6008E284, 32'hDE9178CD);
	test_case(32'hDE684E88, 32'h604AA37F);
	test_case(32'h5FA8B4B6, 32'h60105B29);
	test_case(32'h5FF1EF75, 32'hE04B8381);
	test_case(32'h5F92F4AF, 32'h601035A3);
	test_case(32'hDFE01465, 32'hE0672A78);
	test_case(32'h604BEE64, 32'h604BD288);
	test_case(32'h5F65DFFE, 32'h5FF0B918);
	test_case(32'hDDA179B9, 32'hE0294F67);
	test_case(32'h5FAE5403, 32'hDF1689BA);
	test_case(32'h6030C97C, 32'h5FDA88FA);
	test_case(32'hE065D993, 32'h601C1448);
	test_case(32'hE03F81DA, 32'hE0392E42);
	test_case(32'h5FC0D072, 32'hE077B13C);
	test_case(32'hE077E8A6, 32'h603EDAB0);
	test_case(32'hE070EADC, 32'h604935A4);
	test_case(32'hDF088912, 32'h6043D7FB);
	test_case(32'h5F10574B, 32'h5F5FB3ED);
	test_case(32'h6071D3D5, 32'h5E954C29);
	test_case(32'h5FDFD2F0, 32'hE0575509);
	test_case(32'hDF7E25D3, 32'h6051EFEF);
	test_case(32'h60710134, 32'hE02292CC);
	test_case(32'h60024CD2, 32'hE00358A4);
	test_case(32'h5FE25DBD, 32'h6034D82F);
	test_case(32'h5FB03F3F, 32'h601803EE);
	test_case(32'h604BB975, 32'h5F3225C9);
	test_case(32'h603F7D79, 32'hE06B5566);
	test_case(32'hDFCB3D29, 32'hE05268AB);
	test_case(32'hE0205E22, 32'h60703BFB);
	test_case(32'hE07BB993, 32'h5FD9B358);
	test_case(32'h5DBDF7F4, 32'h607354F9);
	test_case(32'hDF9A2A7F, 32'hE017E25E);
	test_case(32'h5FA4F9BC, 32'h5ED8D47F);
	test_case(32'hE0542CF1, 32'h606A210C);
	test_case(32'h601768B3, 32'hE0130CD6);
	test_case(32'hDFDBD6B7, 32'hDFACDF52);
	test_case(32'h60788192, 32'h602D0542);
	test_case(32'h6024C9C2, 32'h5FCFFF2F);
	test_case(32'h603DAE88, 32'hE04E99D0);
	test_case(32'h604215F9, 32'hE03C8D9C);
	test_case(32'hDD8475E2, 32'hDFA06BA9);
	test_case(32'hE0078B73, 32'hE0081B6D);
	test_case(32'hDED1409E, 32'h5FFAAD2E);
	test_case(32'h600CB7A2, 32'hDF88A8A6);
	test_case(32'hDF032FD8, 32'h5FBADC61);
	test_case(32'h60678C72, 32'hE001F339);
	test_case(32'h5E9E7959, 32'hE01CEB84);
	test_case(32'hE071237D, 32'h6068DD27);
	test_case(32'hDF269241, 32'hDCB84562);
	test_case(32'hE0099C40, 32'h5FFBF732);
	test_case(32'h606086D0, 32'h606465A5);
	test_case(32'hE063BE5C, 32'hDF17CF6A);
	test_case(32'h5FE4B3AC, 32'h604868B5);
	test_case(32'hE041A5A1, 32'h6038A088);
	test_case(32'h5EFAFF9A, 32'hE07057FB);
	test_case(32'hE07B935F, 32'hE05026D4);
	test_case(32'h6013A0BE, 32'hDFE130E7);
	test_case(32'hDF4D48A5, 32'hE03CB22B);
	test_case(32'hDFF69B74, 32'h5FBBF4E6);
	test_case(32'h604676C2, 32'h5FB08F47);
	test_case(32'h607AA309, 32'hE06AC589);
	test_case(32'h5F9E8E6F, 32'hDFC50321);
	test_case(32'h607F0164, 32'h5F93FD91);
	test_case(32'h5FFBDC04, 32'hDF384217);
	test_case(32'h602616FF, 32'h5E6B2718);
	test_case(32'hE00C597B, 32'h60738BF7);
	test_case(32'h5FF51F90, 32'hE002136A);
	test_case(32'h5E1FD44E, 32'h5F39602E);
	test_case(32'h6030D710, 32'hDF8E091F);
	test_case(32'h5F47FBBA, 32'h605B636C);
	test_case(32'h605A965E, 32'h601531E1);
	test_case(32'hDF82920B, 32'hE044F5F9);
	test_case(32'h5FE1CFF4, 32'h603F5FEE);
	test_case(32'h6013C263, 32'h605E8857);
	test_case(32'hDF2927EA, 32'h6072F8F3);
	test_case(32'hE0069884, 32'hDE76F460);
	test_case(32'h5FC2801C, 32'h606CEC5D);
	test_case(32'h60776D21, 32'hE00CB40C);
	test_case(32'h600675C8, 32'h604C2BCD);
	test_case(32'h5FDDBF3B, 32'h5EC38D85);
	test_case(32'h5F9EA04B, 32'h606E4027);
	test_case(32'h605C2BDC, 32'h60319EC8);
	test_case(32'hDFE42711, 32'h5F9C4790);
	test_case(32'hDE9E7300, 32'h601AC083);
	test_case(32'h6042ABD9, 32'h60248A51);
	test_case(32'h5FCCB2D5, 32'h5E2C20A2);
	test_case(32'hDF974E59, 32'hE029E735);
	test_case(32'hE07ABD83, 32'h6011EA61);
	test_case(32'hDFB30BA9, 32'h600FB459);
	test_case(32'h6059D44A, 32'h6017A76B);
	test_case(32'h607C0A74, 32'h5DC88DE1);
	test_case(32'hDF3D938A, 32'hDFC7577B);
	test_case(32'h603B0196, 32'hE070F624);
	test_case(32'hE044A011, 32'h607DD369);
	test_case(32'hDE87B539, 32'hE022DC1B);
	test_case(32'h602EA5DA, 32'h6032D8D7);
	test_case(32'h5FFF540A, 32'hDF2C00FD);
	test_case(32'hE0295B61, 32'h60197134);
	test_case(32'hDFD14B90, 32'hE01B1866);
	test_case(32'h5FC5E226, 32'h5F342BC0);
	test_case(32'h60340F7C, 32'hE0411D78);
	test_case(32'hE059D961, 32'hDFBD39EB);
	test_case(32'h5F93EF17, 32'hDFFAA3CA);
	test_case(32'hDEE8AAE6, 32'h6019C9A8);
	test_case(32'h601ACB3A, 32'h601B521F);
	test_case(32'h5FEABAC9, 32'hE04969F5);
	test_case(32'h600D42FB, 32'hDFB6DA36);
	test_case(32'hDF82BB51, 32'h6000143A);
	test_case(32'h5FE32795, 32'hE025CD63);
	test_case(32'h607FA3F4, 32'h607DAD67);
	test_case(32'hE022EFF4, 32'hDEA3355B);
	test_case(32'h5F8835A7, 32'h5F26195C);
	test_case(32'h607CC232, 32'hDF4BE463);
	test_case(32'h606541D8, 32'hE06DC58E);
	test_case(32'hE0545845, 32'h603FE0A2);
	test_case(32'hE0766F85, 32'hE07ABB54);
	test_case(32'h6016A353, 32'h5FE496BB);
	test_case(32'h5F692ADD, 32'h6007DBCD);
	test_case(32'hDF36EF96, 32'hDF7276BE);
	test_case(32'h5EFE4EBA, 32'h5FC60AD7);
	test_case(32'h6067B0E5, 32'h5F79CF7E);
	test_case(32'hE0231787, 32'h60112666);
	test_case(32'hDF642FB2, 32'h6051E64E);
	test_case(32'h5FB44C41, 32'h5EE2277C);
	test_case(32'h6058C27A, 32'hDF4A01B9);
	test_case(32'hDF811AFC, 32'h60541029);
	test_case(32'h5FEB11D2, 32'hE04128FD);
	test_case(32'h60559043, 32'hDFFCAAF3);
	test_case(32'hDE6E38FF, 32'hDFF99F9A);
	test_case(32'h5F1C5A26, 32'hE046795E);
	test_case(32'h60341878, 32'h5F152276);
	test_case(32'hDE18F235, 32'hDFEAF5E0);
	test_case(32'hDEB5F36E, 32'h5EEF3D0A);
	test_case(32'hE0423059, 32'hE04215AC);
	test_case(32'hE05CB65A, 32'hE073C1AB);
	test_case(32'h6074021E, 32'h5F4B5996);
	test_case(32'hE02B8F7C, 32'h6028359D);
	test_case(32'h6041858E, 32'hE057196C);
	test_case(32'h5F8A956F, 32'hDFA1E3BD);
	test_case(32'h60386632, 32'h605A705B);
	test_case(32'hDF9F5946, 32'hDF999A24);
	test_case(32'h5E1D2B4E, 32'h6068A4F1);
	test_case(32'hDFD96D1A, 32'hE0119542);
	test_case(32'hDF3AAE64, 32'h5FF25DEF);
	test_case(32'h5F8F11C2, 32'hDFDFFBDF);
	test_case(32'hDBA00142, 32'h6011E556);
	test_case(32'h5FC0F51F, 32'hE01B4728);
	test_case(32'h5E7821C6, 32'h5F8DBC1D);
	test_case(32'h5F2338B9, 32'hE07C8036);
	test_case(32'hDE2835DE, 32'hE03287F2);
	test_case(32'hDFBC6220, 32'hDFEBAC01);
	test_case(32'h5FB3D632, 32'h60542B98);
	test_case(32'hE06FC475, 32'hE047E810);
	test_case(32'h5F18859A, 32'hE0505A2E);
	test_case(32'hE015F212, 32'h5DA14ED3);
	test_case(32'h5FE27C2E, 32'hDD69D6BB);
	test_case(32'hE0314489, 32'h5F23EF2C);
	test_case(32'h6030528C, 32'h5E18FA00);
	test_case(32'h607F224E, 32'h6056C350);
	test_case(32'hE01A8CB6, 32'h5F97580D);
	test_case(32'h5F5F511E, 32'hE00FCE97);
	test_case(32'hDF2C7F13, 32'hDF6CE37D);
	test_case(32'h601E396B, 32'hDFB2A383);
	test_case(32'h60798C6C, 32'hDEF18D22);
	test_case(32'hDFE00E20, 32'h5F97934C);
	test_case(32'hE04D60F7, 32'hE04CCB44);
	test_case(32'hDFC1E0DD, 32'hDFDC6099);
	test_case(32'h5FEAFE63, 32'hE05A6FE5);
	test_case(32'h5E8F57C4, 32'h5F9E5E7B);
	test_case(32'hE07D7A5B, 32'h6015B7B0);
	test_case(32'hDF840E7B, 32'h6048816B);
	test_case(32'h60673BEE, 32'hE00956F3);
	test_case(32'hE003063F, 32'hDF400730);
	test_case(32'h5F27E009, 32'h6005F501);
	test_case(32'hE05C81D7, 32'hE05FD25E);
	test_case(32'hDFFF4AF0, 32'hDFD70F1F);
	test_case(32'hE028B0E1, 32'h5FDDD6E2);
	test_case(32'h5F41CEAA, 32'h5F4AF763);
	test_case(32'hE00A786A, 32'h6073D1DB);
	test_case(32'h5F9A9331, 32'h5F47927F);
	test_case(32'hDD6A4FB2, 32'hDF5FB050);
	test_case(32'hE03B21A0, 32'hDE1CAC32);
	test_case(32'hDEDA4F82, 32'h5FEFC27A);
	test_case(32'h5F5BF55F, 32'hDBAD902E);
	test_case(32'hDF58F698, 32'hE0598A84);
	test_case(32'hDF82EFC2, 32'hE0196371);
	test_case(32'h5FB7BCF9, 32'hE03A039A);
	test_case(32'h601BE36F, 32'h5F15F815);
	test_case(32'h5FA2DD64, 32'hDE966ADA);
	test_case(32'h60748C8B, 32'h6040B5AD);
	test_case(32'hDF76C7FB, 32'h5F0AA4BF);
	test_case(32'h5F80CA29, 32'hDF0BB9A2);
	test_case(32'hE04172B8, 32'hDDC7B8AB);
	test_case(32'hE05987AF, 32'h60047596);
	test_case(32'hE05D6459, 32'h605B9DEC);
	test_case(32'h5E8551B3, 32'hE0555D4A);
	test_case(32'hDEDAF277, 32'hDEE3E87E);
	test_case(32'h60789F2D, 32'h60450F1D);
	test_case(32'hDE85CE92, 32'hE02B2529);
	test_case(32'hE03A5E09, 32'h5F75C50F);
	test_case(32'hDF2BBE8B, 32'hDF70E61B);
	test_case(32'h5F00421C, 32'h5FE5EF0B);
	test_case(32'hE03152E5, 32'hE07B5E97);
	test_case(32'hE01C3344, 32'hE06A6C07);
	test_case(32'hDF112029, 32'hDEB03ACA);
	test_case(32'hE01F1919, 32'h5F8D3F60);
	test_case(32'hDEDF204A, 32'hDFB4D519);
	test_case(32'h5E9EC3B9, 32'h604BB1A3);
	test_case(32'hDEC7D6F0, 32'h604E6B34);
	test_case(32'h5CB34420, 32'h6007AF72);
	test_case(32'hE06886F2, 32'hDEBF7D58);
	test_case(32'hDF27912D, 32'hDFF2CDCF);
	test_case(32'hDF27ADA0, 32'h5EA32990);
	test_case(32'hDFD5AA44, 32'hE00E4A2C);
	test_case(32'h5FA9FE03, 32'hDFACA026);
	test_case(32'h5F3468A3, 32'hDF2035D1);
	test_case(32'h60779C03, 32'hDFA30592);
	test_case(32'h601AE12F, 32'h5FF30A1F);
	test_case(32'hDF744984, 32'hE006B1BA);

    $finish;
end

task test_case(
    input [31:0] a_in,
    input [31:0] b_in
); begin
    @(negedge clk) begin
        a = a_in;
        b = b_in;
    end
    @(posedge clk) begin
        $display("%h,%h,%h", a_in, b_in, out);
    end
end
endtask

endmodule
